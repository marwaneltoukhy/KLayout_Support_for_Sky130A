*
*  /home/marwan/ef/klayout_lvs/lvs/test_cases/xres_buf/xres_buf.spice : SPICE netlist translated from the VERILOG netlist : /home/marwan/ef/caravel/verilog/gl/xres_buf.v
*                                                                       on the 2021-12-22 17:58:44.519025
*
***************************************************************************************************************************************************************************

.INCLUDE sky130_fd_sc_hd.spice 

.GLOBAL VDD VSS

.SUBCKT XRES_BUF(A A LVGND LVPWR VGND VPWR X 


.ENDS XRES_BUF(A,