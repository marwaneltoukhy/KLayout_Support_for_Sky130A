*SPICE netlist created from verilog structural netlist module user_id_programming by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /home/marwan/klayout_lvs/lvs/test_cases/user_id_programming/sky130_fd_sc_hd.spice

.subckt user_id_programming VGND VPWR mask_rev[0] mask_rev[1] mask_rev[2] mask_rev[3] mask_rev[4]
+ mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mask_rev[10] mask_rev[11] mask_rev[12]
+ mask_rev[13] mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[20]
+ mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28]
+ mask_rev[29] mask_rev[30] mask_rev[31] 

XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_19 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X\mask_rev_value[0]  VGND VGND VPWR VPWR \user_proj_id_high[0]\ mask_rev[0] sky130_fd_sc_hd__conb_1
X\mask_rev_value[10]  VGND VGND VPWR VPWR \user_proj_id_high[10]\ mask_rev[10] sky130_fd_sc_hd__conb_1
X\mask_rev_value[11]  VGND VGND VPWR VPWR \user_proj_id_high[11]\ mask_rev[11] sky130_fd_sc_hd__conb_1
X\mask_rev_value[12]  VGND VGND VPWR VPWR \user_proj_id_high[12]\ mask_rev[12] sky130_fd_sc_hd__conb_1
X\mask_rev_value[13]  VGND VGND VPWR VPWR \user_proj_id_high[13]\ mask_rev[13] sky130_fd_sc_hd__conb_1
X\mask_rev_value[14]  VGND VGND VPWR VPWR \user_proj_id_high[14]\ mask_rev[14] sky130_fd_sc_hd__conb_1
X\mask_rev_value[15]  VGND VGND VPWR VPWR \user_proj_id_high[15]\ mask_rev[15] sky130_fd_sc_hd__conb_1
X\mask_rev_value[16]  VGND VGND VPWR VPWR \user_proj_id_high[16]\ mask_rev[16] sky130_fd_sc_hd__conb_1
X\mask_rev_value[17]  VGND VGND VPWR VPWR \user_proj_id_high[17]\ mask_rev[17] sky130_fd_sc_hd__conb_1
X\mask_rev_value[18]  VGND VGND VPWR VPWR \user_proj_id_high[18]\ mask_rev[18] sky130_fd_sc_hd__conb_1
X\mask_rev_value[19]  VGND VGND VPWR VPWR \user_proj_id_high[19]\ mask_rev[19] sky130_fd_sc_hd__conb_1
X\mask_rev_value[1]  VGND VGND VPWR VPWR \user_proj_id_high[1]\ mask_rev[1] sky130_fd_sc_hd__conb_1
X\mask_rev_value[20]  VGND VGND VPWR VPWR \user_proj_id_high[20]\ mask_rev[20] sky130_fd_sc_hd__conb_1
X\mask_rev_value[21]  VGND VGND VPWR VPWR \user_proj_id_high[21]\ mask_rev[21] sky130_fd_sc_hd__conb_1
X\mask_rev_value[22]  VGND VGND VPWR VPWR \user_proj_id_high[22]\ mask_rev[22] sky130_fd_sc_hd__conb_1
X\mask_rev_value[23]  VGND VGND VPWR VPWR \user_proj_id_high[23]\ mask_rev[23] sky130_fd_sc_hd__conb_1
X\mask_rev_value[24]  VGND VGND VPWR VPWR \user_proj_id_high[24]\ mask_rev[24] sky130_fd_sc_hd__conb_1
X\mask_rev_value[25]  VGND VGND VPWR VPWR \user_proj_id_high[25]\ mask_rev[25] sky130_fd_sc_hd__conb_1
X\mask_rev_value[26]  VGND VGND VPWR VPWR \user_proj_id_high[26]\ mask_rev[26] sky130_fd_sc_hd__conb_1
X\mask_rev_value[27]  VGND VGND VPWR VPWR \user_proj_id_high[27]\ mask_rev[27] sky130_fd_sc_hd__conb_1
X\mask_rev_value[28]  VGND VGND VPWR VPWR \user_proj_id_high[28]\ mask_rev[28] sky130_fd_sc_hd__conb_1
X\mask_rev_value[29]  VGND VGND VPWR VPWR \user_proj_id_high[29]\ mask_rev[29] sky130_fd_sc_hd__conb_1
X\mask_rev_value[2]  VGND VGND VPWR VPWR \user_proj_id_high[2]\ mask_rev[2] sky130_fd_sc_hd__conb_1
X\mask_rev_value[30]  VGND VGND VPWR VPWR \user_proj_id_high[30]\ mask_rev[30] sky130_fd_sc_hd__conb_1
X\mask_rev_value[31]  VGND VGND VPWR VPWR \user_proj_id_high[31]\ mask_rev[31] sky130_fd_sc_hd__conb_1
X\mask_rev_value[3]  VGND VGND VPWR VPWR \user_proj_id_high[3]\ mask_rev[3] sky130_fd_sc_hd__conb_1
X\mask_rev_value[4]  VGND VGND VPWR VPWR \user_proj_id_high[4]\ mask_rev[4] sky130_fd_sc_hd__conb_1
X\mask_rev_value[5]  VGND VGND VPWR VPWR \user_proj_id_high[5]\ mask_rev[5] sky130_fd_sc_hd__conb_1
X\mask_rev_value[6]  VGND VGND VPWR VPWR \user_proj_id_high[6]\ mask_rev[6] sky130_fd_sc_hd__conb_1
X\mask_rev_value[7]  VGND VGND VPWR VPWR \user_proj_id_high[7]\ mask_rev[7] sky130_fd_sc_hd__conb_1
X\mask_rev_value[8]  VGND VGND VPWR VPWR \user_proj_id_high[8]\ mask_rev[8] sky130_fd_sc_hd__conb_1
X\mask_rev_value[9]  VGND VGND VPWR VPWR \user_proj_id_high[9]\ mask_rev[9] sky130_fd_sc_hd__conb_1

.ends
.end
