*
*  /home/marwan/ef/klayout_lvs/lvs/test_cases/chip_io/chip_io.spice : SPICE netlist translated from the VERILOG netlist : /home/marwan/ef/caravel/verilog/gl/chip_io.v
*                                                                     on the 2021-12-22 17:54:36.053268
*
************************************************************************************************************************************************************************

.INCLUDE sky130_fd_sc_hd.spice 

.GLOBAL VDD VSS

.SUBCKT CHIP_IO(VDDIO_PAD CLOCK CLOCK_CORE FLASH_CLK FLASH_CLK_CORE FLASH_CLK_IEB_CORE FLASH_CLK_OEB_CORE FLASH_CSB FLASH_CSB_CORE FLASH_CSB_IEB_CORE FLASH_CSB_OEB_CORE FLASH_IO0 FLASH_IO0_DI_CORE FLASH_IO0_DO_CORE FLASH_IO0_IEB_CORE FLASH_IO0_OEB_CORE FLASH_IO1 FLASH_IO1_DI_CORE FLASH_IO1_DO_CORE FLASH_IO1_IEB_CORE FLASH_IO1_OEB_CORE GPIO GPIO_IN_CORE GPIO_INENB_CORE GPIO_MODE0_CORE GPIO_MODE1_CORE GPIO_OUT_CORE GPIO_OUTENB_CORE MPRJ_ANALOG_IO[0] MPRJ_ANALOG_IO[1] MPRJ_ANALOG_IO[2] MPRJ_ANALOG_IO[3] MPRJ_ANALOG_IO[4] MPRJ_ANALOG_IO[5] MPRJ_ANALOG_IO[6] MPRJ_ANALOG_IO[7] MPRJ_ANALOG_IO[8] MPRJ_ANALOG_IO[9] MPRJ_ANALOG_IO[10] MPRJ_ANALOG_IO[11] MPRJ_ANALOG_IO[12] MPRJ_ANALOG_IO[13] MPRJ_ANALOG_IO[14] MPRJ_ANALOG_IO[15] MPRJ_ANALOG_IO[16] MPRJ_ANALOG_IO[17] MPRJ_ANALOG_IO[18] MPRJ_ANALOG_IO[19] MPRJ_ANALOG_IO[20] MPRJ_ANALOG_IO[21] MPRJ_ANALOG_IO[22] MPRJ_ANALOG_IO[23] MPRJ_ANALOG_IO[24] MPRJ_ANALOG_IO[25] MPRJ_ANALOG_IO[26] MPRJ_ANALOG_IO[27] MPRJ_ANALOG_IO[28] MPRJ_IO[0] MPRJ_IO[1] MPRJ_IO[2] MPRJ_IO[3] MPRJ_IO[4] MPRJ_IO[5] MPRJ_IO[6] MPRJ_IO[7] MPRJ_IO[8] MPRJ_IO[9] MPRJ_IO[10] MPRJ_IO[11] MPRJ_IO[12] MPRJ_IO[13] MPRJ_IO[14] MPRJ_IO[15] MPRJ_IO[16] MPRJ_IO[17] MPRJ_IO[18] MPRJ_IO[19] MPRJ_IO[20] MPRJ_IO[21] MPRJ_IO[22] MPRJ_IO[23] MPRJ_IO[24] MPRJ_IO[25] MPRJ_IO[26] MPRJ_IO[27] MPRJ_IO[28] MPRJ_IO[29] MPRJ_IO[30] MPRJ_IO[31] MPRJ_IO[32] MPRJ_IO[33] MPRJ_IO[34] MPRJ_IO[35] MPRJ_IO[36] MPRJ_IO[37] MPRJ_IO_ANALOG_EN[0] MPRJ_IO_ANALOG_EN[1] MPRJ_IO_ANALOG_EN[2] MPRJ_IO_ANALOG_EN[3] MPRJ_IO_ANALOG_EN[4] MPRJ_IO_ANALOG_EN[5] MPRJ_IO_ANALOG_EN[6] MPRJ_IO_ANALOG_EN[7] MPRJ_IO_ANALOG_EN[8] MPRJ_IO_ANALOG_EN[9] MPRJ_IO_ANALOG_EN[10] MPRJ_IO_ANALOG_EN[11] MPRJ_IO_ANALOG_EN[12] MPRJ_IO_ANALOG_EN[13] MPRJ_IO_ANALOG_EN[14] MPRJ_IO_ANALOG_EN[15] MPRJ_IO_ANALOG_EN[16] MPRJ_IO_ANALOG_EN[17] MPRJ_IO_ANALOG_EN[18] MPRJ_IO_ANALOG_EN[19] MPRJ_IO_ANALOG_EN[20] MPRJ_IO_ANALOG_EN[21] MPRJ_IO_ANALOG_EN[22] MPRJ_IO_ANALOG_EN[23] MPRJ_IO_ANALOG_EN[24] MPRJ_IO_ANALOG_EN[25] MPRJ_IO_ANALOG_EN[26] MPRJ_IO_ANALOG_EN[27] MPRJ_IO_ANALOG_EN[28] MPRJ_IO_ANALOG_EN[29] MPRJ_IO_ANALOG_EN[30] MPRJ_IO_ANALOG_EN[31] MPRJ_IO_ANALOG_EN[32] MPRJ_IO_ANALOG_EN[33] MPRJ_IO_ANALOG_EN[34] MPRJ_IO_ANALOG_EN[35] MPRJ_IO_ANALOG_EN[36] MPRJ_IO_ANALOG_EN[37] MPRJ_IO_ANALOG_POL[0] MPRJ_IO_ANALOG_POL[1] MPRJ_IO_ANALOG_POL[2] MPRJ_IO_ANALOG_POL[3] MPRJ_IO_ANALOG_POL[4] MPRJ_IO_ANALOG_POL[5] MPRJ_IO_ANALOG_POL[6] MPRJ_IO_ANALOG_POL[7] MPRJ_IO_ANALOG_POL[8] MPRJ_IO_ANALOG_POL[9] MPRJ_IO_ANALOG_POL[10] MPRJ_IO_ANALOG_POL[11] MPRJ_IO_ANALOG_POL[12] MPRJ_IO_ANALOG_POL[13] MPRJ_IO_ANALOG_POL[14] MPRJ_IO_ANALOG_POL[15] MPRJ_IO_ANALOG_POL[16] MPRJ_IO_ANALOG_POL[17] MPRJ_IO_ANALOG_POL[18] MPRJ_IO_ANALOG_POL[19] MPRJ_IO_ANALOG_POL[20] MPRJ_IO_ANALOG_POL[21] MPRJ_IO_ANALOG_POL[22] MPRJ_IO_ANALOG_POL[23] MPRJ_IO_ANALOG_POL[24] MPRJ_IO_ANALOG_POL[25] MPRJ_IO_ANALOG_POL[26] MPRJ_IO_ANALOG_POL[27] MPRJ_IO_ANALOG_POL[28] MPRJ_IO_ANALOG_POL[29] MPRJ_IO_ANALOG_POL[30] MPRJ_IO_ANALOG_POL[31] MPRJ_IO_ANALOG_POL[32] MPRJ_IO_ANALOG_POL[33] MPRJ_IO_ANALOG_POL[34] MPRJ_IO_ANALOG_POL[35] MPRJ_IO_ANALOG_POL[36] MPRJ_IO_ANALOG_POL[37] MPRJ_IO_ANALOG_SEL[0] MPRJ_IO_ANALOG_SEL[1] MPRJ_IO_ANALOG_SEL[2] MPRJ_IO_ANALOG_SEL[3] MPRJ_IO_ANALOG_SEL[4] MPRJ_IO_ANALOG_SEL[5] MPRJ_IO_ANALOG_SEL[6] MPRJ_IO_ANALOG_SEL[7] MPRJ_IO_ANALOG_SEL[8] MPRJ_IO_ANALOG_SEL[9] MPRJ_IO_ANALOG_SEL[10] MPRJ_IO_ANALOG_SEL[11] MPRJ_IO_ANALOG_SEL[12] MPRJ_IO_ANALOG_SEL[13] MPRJ_IO_ANALOG_SEL[14] MPRJ_IO_ANALOG_SEL[15] MPRJ_IO_ANALOG_SEL[16] MPRJ_IO_ANALOG_SEL[17] MPRJ_IO_ANALOG_SEL[18] MPRJ_IO_ANALOG_SEL[19] MPRJ_IO_ANALOG_SEL[20] MPRJ_IO_ANALOG_SEL[21] MPRJ_IO_ANALOG_SEL[22] MPRJ_IO_ANALOG_SEL[23] MPRJ_IO_ANALOG_SEL[24] MPRJ_IO_ANALOG_SEL[25] MPRJ_IO_ANALOG_SEL[26] MPRJ_IO_ANALOG_SEL[27] MPRJ_IO_ANALOG_SEL[28] MPRJ_IO_ANALOG_SEL[29] MPRJ_IO_ANALOG_SEL[30] MPRJ_IO_ANALOG_SEL[31] MPRJ_IO_ANALOG_SEL[32] MPRJ_IO_ANALOG_SEL[33] MPRJ_IO_ANALOG_SEL[34] MPRJ_IO_ANALOG_SEL[35] MPRJ_IO_ANALOG_SEL[36] MPRJ_IO_ANALOG_SEL[37] MPRJ_IO_DM[0] MPRJ_IO_DM[1] MPRJ_IO_DM[2] MPRJ_IO_DM[3] MPRJ_IO_DM[4] MPRJ_IO_DM[5] MPRJ_IO_DM[6] MPRJ_IO_DM[7] MPRJ_IO_DM[8] MPRJ_IO_DM[9] MPRJ_IO_DM[10] MPRJ_IO_DM[11] MPRJ_IO_DM[12] MPRJ_IO_DM[13] MPRJ_IO_DM[14] MPRJ_IO_DM[15] MPRJ_IO_DM[16] MPRJ_IO_DM[17] MPRJ_IO_DM[18] MPRJ_IO_DM[19] MPRJ_IO_DM[20] MPRJ_IO_DM[21] MPRJ_IO_DM[22] MPRJ_IO_DM[23] MPRJ_IO_DM[24] MPRJ_IO_DM[25] MPRJ_IO_DM[26] MPRJ_IO_DM[27] MPRJ_IO_DM[28] MPRJ_IO_DM[29] MPRJ_IO_DM[30] MPRJ_IO_DM[31] MPRJ_IO_DM[32] MPRJ_IO_DM[33] MPRJ_IO_DM[34] MPRJ_IO_DM[35] MPRJ_IO_DM[36] MPRJ_IO_DM[37] MPRJ_IO_DM[38] MPRJ_IO_DM[39] MPRJ_IO_DM[40] MPRJ_IO_DM[41] MPRJ_IO_DM[42] MPRJ_IO_DM[43] MPRJ_IO_DM[44] MPRJ_IO_DM[45] MPRJ_IO_DM[46] MPRJ_IO_DM[47] MPRJ_IO_DM[48] MPRJ_IO_DM[49] MPRJ_IO_DM[50] MPRJ_IO_DM[51] MPRJ_IO_DM[52] MPRJ_IO_DM[53] MPRJ_IO_DM[54] MPRJ_IO_DM[55] MPRJ_IO_DM[56] MPRJ_IO_DM[57] MPRJ_IO_DM[58] MPRJ_IO_DM[59] MPRJ_IO_DM[60] MPRJ_IO_DM[61] MPRJ_IO_DM[62] MPRJ_IO_DM[63] MPRJ_IO_DM[64] MPRJ_IO_DM[65] MPRJ_IO_DM[66] MPRJ_IO_DM[67] MPRJ_IO_DM[68] MPRJ_IO_DM[69] MPRJ_IO_DM[70] MPRJ_IO_DM[71] MPRJ_IO_DM[72] MPRJ_IO_DM[73] MPRJ_IO_DM[74] MPRJ_IO_DM[75] MPRJ_IO_DM[76] MPRJ_IO_DM[77] MPRJ_IO_DM[78] MPRJ_IO_DM[79] MPRJ_IO_DM[80] MPRJ_IO_DM[81] MPRJ_IO_DM[82] MPRJ_IO_DM[83] MPRJ_IO_DM[84] MPRJ_IO_DM[85] MPRJ_IO_DM[86] MPRJ_IO_DM[87] MPRJ_IO_DM[88] MPRJ_IO_DM[89] MPRJ_IO_DM[90] MPRJ_IO_DM[91] MPRJ_IO_DM[92] MPRJ_IO_DM[93] MPRJ_IO_DM[94] MPRJ_IO_DM[95] MPRJ_IO_DM[96] MPRJ_IO_DM[97] MPRJ_IO_DM[98] MPRJ_IO_DM[99] MPRJ_IO_DM[100] MPRJ_IO_DM[101] MPRJ_IO_DM[102] MPRJ_IO_DM[103] MPRJ_IO_DM[104] MPRJ_IO_DM[105] MPRJ_IO_DM[106] MPRJ_IO_DM[107] MPRJ_IO_DM[108] MPRJ_IO_DM[109] MPRJ_IO_DM[110] MPRJ_IO_DM[111] MPRJ_IO_DM[112] MPRJ_IO_DM[113] MPRJ_IO_HOLDOVER[0] MPRJ_IO_HOLDOVER[1] MPRJ_IO_HOLDOVER[2] MPRJ_IO_HOLDOVER[3] MPRJ_IO_HOLDOVER[4] MPRJ_IO_HOLDOVER[5] MPRJ_IO_HOLDOVER[6] MPRJ_IO_HOLDOVER[7] MPRJ_IO_HOLDOVER[8] MPRJ_IO_HOLDOVER[9] MPRJ_IO_HOLDOVER[10] MPRJ_IO_HOLDOVER[11] MPRJ_IO_HOLDOVER[12] MPRJ_IO_HOLDOVER[13] MPRJ_IO_HOLDOVER[14] MPRJ_IO_HOLDOVER[15] MPRJ_IO_HOLDOVER[16] MPRJ_IO_HOLDOVER[17] MPRJ_IO_HOLDOVER[18] MPRJ_IO_HOLDOVER[19] MPRJ_IO_HOLDOVER[20] MPRJ_IO_HOLDOVER[21] MPRJ_IO_HOLDOVER[22] MPRJ_IO_HOLDOVER[23] MPRJ_IO_HOLDOVER[24] MPRJ_IO_HOLDOVER[25] MPRJ_IO_HOLDOVER[26] MPRJ_IO_HOLDOVER[27] MPRJ_IO_HOLDOVER[28] MPRJ_IO_HOLDOVER[29] MPRJ_IO_HOLDOVER[30] MPRJ_IO_HOLDOVER[31] MPRJ_IO_HOLDOVER[32] MPRJ_IO_HOLDOVER[33] MPRJ_IO_HOLDOVER[34] MPRJ_IO_HOLDOVER[35] MPRJ_IO_HOLDOVER[36] MPRJ_IO_HOLDOVER[37] MPRJ_IO_IB_MODE_SEL[0] MPRJ_IO_IB_MODE_SEL[1] MPRJ_IO_IB_MODE_SEL[2] MPRJ_IO_IB_MODE_SEL[3] MPRJ_IO_IB_MODE_SEL[4] MPRJ_IO_IB_MODE_SEL[5] MPRJ_IO_IB_MODE_SEL[6] MPRJ_IO_IB_MODE_SEL[7] MPRJ_IO_IB_MODE_SEL[8] MPRJ_IO_IB_MODE_SEL[9] MPRJ_IO_IB_MODE_SEL[10] MPRJ_IO_IB_MODE_SEL[11] MPRJ_IO_IB_MODE_SEL[12] MPRJ_IO_IB_MODE_SEL[13] MPRJ_IO_IB_MODE_SEL[14] MPRJ_IO_IB_MODE_SEL[15] MPRJ_IO_IB_MODE_SEL[16] MPRJ_IO_IB_MODE_SEL[17] MPRJ_IO_IB_MODE_SEL[18] MPRJ_IO_IB_MODE_SEL[19] MPRJ_IO_IB_MODE_SEL[20] MPRJ_IO_IB_MODE_SEL[21] MPRJ_IO_IB_MODE_SEL[22] MPRJ_IO_IB_MODE_SEL[23] MPRJ_IO_IB_MODE_SEL[24] MPRJ_IO_IB_MODE_SEL[25] MPRJ_IO_IB_MODE_SEL[26] MPRJ_IO_IB_MODE_SEL[27] MPRJ_IO_IB_MODE_SEL[28] MPRJ_IO_IB_MODE_SEL[29] MPRJ_IO_IB_MODE_SEL[30] MPRJ_IO_IB_MODE_SEL[31] MPRJ_IO_IB_MODE_SEL[32] MPRJ_IO_IB_MODE_SEL[33] MPRJ_IO_IB_MODE_SEL[34] MPRJ_IO_IB_MODE_SEL[35] MPRJ_IO_IB_MODE_SEL[36] MPRJ_IO_IB_MODE_SEL[37] MPRJ_IO_IN[0] MPRJ_IO_IN[1] MPRJ_IO_IN[2] MPRJ_IO_IN[3] MPRJ_IO_IN[4] MPRJ_IO_IN[5] MPRJ_IO_IN[6] MPRJ_IO_IN[7] MPRJ_IO_IN[8] MPRJ_IO_IN[9] MPRJ_IO_IN[10] MPRJ_IO_IN[11] MPRJ_IO_IN[12] MPRJ_IO_IN[13] MPRJ_IO_IN[14] MPRJ_IO_IN[15] MPRJ_IO_IN[16] MPRJ_IO_IN[17] MPRJ_IO_IN[18] MPRJ_IO_IN[19] MPRJ_IO_IN[20] MPRJ_IO_IN[21] MPRJ_IO_IN[22] MPRJ_IO_IN[23] MPRJ_IO_IN[24] MPRJ_IO_IN[25] MPRJ_IO_IN[26] MPRJ_IO_IN[27] MPRJ_IO_IN[28] MPRJ_IO_IN[29] MPRJ_IO_IN[30] MPRJ_IO_IN[31] MPRJ_IO_IN[32] MPRJ_IO_IN[33] MPRJ_IO_IN[34] MPRJ_IO_IN[35] MPRJ_IO_IN[36] MPRJ_IO_IN[37] MPRJ_IO_INP_DIS[0] MPRJ_IO_INP_DIS[1] MPRJ_IO_INP_DIS[2] MPRJ_IO_INP_DIS[3] MPRJ_IO_INP_DIS[4] MPRJ_IO_INP_DIS[5] MPRJ_IO_INP_DIS[6] MPRJ_IO_INP_DIS[7] MPRJ_IO_INP_DIS[8] MPRJ_IO_INP_DIS[9] MPRJ_IO_INP_DIS[10] MPRJ_IO_INP_DIS[11] MPRJ_IO_INP_DIS[12] MPRJ_IO_INP_DIS[13] MPRJ_IO_INP_DIS[14] MPRJ_IO_INP_DIS[15] MPRJ_IO_INP_DIS[16] MPRJ_IO_INP_DIS[17] MPRJ_IO_INP_DIS[18] MPRJ_IO_INP_DIS[19] MPRJ_IO_INP_DIS[20] MPRJ_IO_INP_DIS[21] MPRJ_IO_INP_DIS[22] MPRJ_IO_INP_DIS[23] MPRJ_IO_INP_DIS[24] MPRJ_IO_INP_DIS[25] MPRJ_IO_INP_DIS[26] MPRJ_IO_INP_DIS[27] MPRJ_IO_INP_DIS[28] MPRJ_IO_INP_DIS[29] MPRJ_IO_INP_DIS[30] MPRJ_IO_INP_DIS[31] MPRJ_IO_INP_DIS[32] MPRJ_IO_INP_DIS[33] MPRJ_IO_INP_DIS[34] MPRJ_IO_INP_DIS[35] MPRJ_IO_INP_DIS[36] MPRJ_IO_INP_DIS[37] MPRJ_IO_OEB[0] MPRJ_IO_OEB[1] MPRJ_IO_OEB[2] MPRJ_IO_OEB[3] MPRJ_IO_OEB[4] MPRJ_IO_OEB[5] MPRJ_IO_OEB[6] MPRJ_IO_OEB[7] MPRJ_IO_OEB[8] MPRJ_IO_OEB[9] MPRJ_IO_OEB[10] MPRJ_IO_OEB[11] MPRJ_IO_OEB[12] MPRJ_IO_OEB[13] MPRJ_IO_OEB[14] MPRJ_IO_OEB[15] MPRJ_IO_OEB[16] MPRJ_IO_OEB[17] MPRJ_IO_OEB[18] MPRJ_IO_OEB[19] MPRJ_IO_OEB[20] MPRJ_IO_OEB[21] MPRJ_IO_OEB[22] MPRJ_IO_OEB[23] MPRJ_IO_OEB[24] MPRJ_IO_OEB[25] MPRJ_IO_OEB[26] MPRJ_IO_OEB[27] MPRJ_IO_OEB[28] MPRJ_IO_OEB[29] MPRJ_IO_OEB[30] MPRJ_IO_OEB[31] MPRJ_IO_OEB[32] MPRJ_IO_OEB[33] MPRJ_IO_OEB[34] MPRJ_IO_OEB[35] MPRJ_IO_OEB[36] MPRJ_IO_OEB[37] MPRJ_IO_OUT[0] MPRJ_IO_OUT[1] MPRJ_IO_OUT[2] MPRJ_IO_OUT[3] MPRJ_IO_OUT[4] MPRJ_IO_OUT[5] MPRJ_IO_OUT[6] MPRJ_IO_OUT[7] MPRJ_IO_OUT[8] MPRJ_IO_OUT[9] MPRJ_IO_OUT[10] MPRJ_IO_OUT[11] MPRJ_IO_OUT[12] MPRJ_IO_OUT[13] MPRJ_IO_OUT[14] MPRJ_IO_OUT[15] MPRJ_IO_OUT[16] MPRJ_IO_OUT[17] MPRJ_IO_OUT[18] MPRJ_IO_OUT[19] MPRJ_IO_OUT[20] MPRJ_IO_OUT[21] MPRJ_IO_OUT[22] MPRJ_IO_OUT[23] MPRJ_IO_OUT[24] MPRJ_IO_OUT[25] MPRJ_IO_OUT[26] MPRJ_IO_OUT[27] MPRJ_IO_OUT[28] MPRJ_IO_OUT[29] MPRJ_IO_OUT[30] MPRJ_IO_OUT[31] MPRJ_IO_OUT[32] MPRJ_IO_OUT[33] MPRJ_IO_OUT[34] MPRJ_IO_OUT[35] MPRJ_IO_OUT[36] MPRJ_IO_OUT[37] MPRJ_IO_SLOW_SEL[0] MPRJ_IO_SLOW_SEL[1] MPRJ_IO_SLOW_SEL[2] MPRJ_IO_SLOW_SEL[3] MPRJ_IO_SLOW_SEL[4] MPRJ_IO_SLOW_SEL[5] MPRJ_IO_SLOW_SEL[6] MPRJ_IO_SLOW_SEL[7] MPRJ_IO_SLOW_SEL[8] MPRJ_IO_SLOW_SEL[9] MPRJ_IO_SLOW_SEL[10] MPRJ_IO_SLOW_SEL[11] MPRJ_IO_SLOW_SEL[12] MPRJ_IO_SLOW_SEL[13] MPRJ_IO_SLOW_SEL[14] MPRJ_IO_SLOW_SEL[15] MPRJ_IO_SLOW_SEL[16] MPRJ_IO_SLOW_SEL[17] MPRJ_IO_SLOW_SEL[18] MPRJ_IO_SLOW_SEL[19] MPRJ_IO_SLOW_SEL[20] MPRJ_IO_SLOW_SEL[21] MPRJ_IO_SLOW_SEL[22] MPRJ_IO_SLOW_SEL[23] MPRJ_IO_SLOW_SEL[24] MPRJ_IO_SLOW_SEL[25] MPRJ_IO_SLOW_SEL[26] MPRJ_IO_SLOW_SEL[27] MPRJ_IO_SLOW_SEL[28] MPRJ_IO_SLOW_SEL[29] MPRJ_IO_SLOW_SEL[30] MPRJ_IO_SLOW_SEL[31] MPRJ_IO_SLOW_SEL[32] MPRJ_IO_SLOW_SEL[33] MPRJ_IO_SLOW_SEL[34] MPRJ_IO_SLOW_SEL[35] MPRJ_IO_SLOW_SEL[36] MPRJ_IO_SLOW_SEL[37] MPRJ_IO_VTRIP_SEL[0] MPRJ_IO_VTRIP_SEL[1] MPRJ_IO_VTRIP_SEL[2] MPRJ_IO_VTRIP_SEL[3] MPRJ_IO_VTRIP_SEL[4] MPRJ_IO_VTRIP_SEL[5] MPRJ_IO_VTRIP_SEL[6] MPRJ_IO_VTRIP_SEL[7] MPRJ_IO_VTRIP_SEL[8] MPRJ_IO_VTRIP_SEL[9] MPRJ_IO_VTRIP_SEL[10] MPRJ_IO_VTRIP_SEL[11] MPRJ_IO_VTRIP_SEL[12] MPRJ_IO_VTRIP_SEL[13] MPRJ_IO_VTRIP_SEL[14] MPRJ_IO_VTRIP_SEL[15] MPRJ_IO_VTRIP_SEL[16] MPRJ_IO_VTRIP_SEL[17] MPRJ_IO_VTRIP_SEL[18] MPRJ_IO_VTRIP_SEL[19] MPRJ_IO_VTRIP_SEL[20] MPRJ_IO_VTRIP_SEL[21] MPRJ_IO_VTRIP_SEL[22] MPRJ_IO_VTRIP_SEL[23] MPRJ_IO_VTRIP_SEL[24] MPRJ_IO_VTRIP_SEL[25] MPRJ_IO_VTRIP_SEL[26] MPRJ_IO_VTRIP_SEL[27] MPRJ_IO_VTRIP_SEL[28] MPRJ_IO_VTRIP_SEL[29] MPRJ_IO_VTRIP_SEL[30] MPRJ_IO_VTRIP_SEL[31] MPRJ_IO_VTRIP_SEL[32] MPRJ_IO_VTRIP_SEL[33] MPRJ_IO_VTRIP_SEL[34] MPRJ_IO_VTRIP_SEL[35] MPRJ_IO_VTRIP_SEL[36] MPRJ_IO_VTRIP_SEL[37] POR PORB_H RESETB RESETB_CORE_H VCCD VCCD1 VCCD1_PAD VCCD2 VCCD2_PAD VCCD_PAD VDDA VDDA1 VDDA1_PAD VDDA1_PAD2 VDDA2 VDDA2_PAD VDDA_PAD VDDIO VDDIO_PAD VDDIO_PAD2 VSSA VSSA1 VSSA1_PAD VSSA1_PAD2 VSSA2 VSSA2_PAD VSSA_PAD VSSD VSSD1 VSSD1_PAD VSSD2 VSSD2_PAD VSSD_PAD VSSIO VSSIO_PAD VSSIO_PAD2 


.ENDS CHIP_IO(VDDIO_PAD,