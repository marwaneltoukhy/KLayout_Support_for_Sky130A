* Extracted by KLayout on : 19/01/2022 09:20

.SUBCKT housekeeping pad_flash_clk_oeb pad_flash_csb pad_flash_csb_oeb
+ pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb pad_flash_io0_oeb
+ pad_flash_io1_di pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb
+ pll_dco_ena pll_div[0] pll_div[1] pll_div[2] pll_div[3] pll_div[4] pll_sel[0]
+ pll_sel[1] pll_sel[2] pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_trim[0]
+ pll_trim[1] pll_trim[2] pll_trim[3] pll_trim[4] pll_trim[5] pll_trim[6]
+ pll_trim[7] pll_trim[8] pll_trim[9] pll_trim[10] pll_trim[11] pll_trim[12]
+ pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16] pll_trim[17] pll_trim[18]
+ pll_trim[19] pll_trim[20] pll_trim[21] pll_trim[22] pll_trim[23] pll_trim[24]
+ pll_trim[25] pll_bypass mask_rev_in[0] mask_rev_in[1] mask_rev_in[2]
+ mask_rev_in[3] mask_rev_in[4] mask_rev_in[5] mask_rev_in[6] mask_rev_in[7]
+ mask_rev_in[8] mask_rev_in[9] mask_rev_in[10] mask_rev_in[11] mask_rev_in[12]
+ mask_rev_in[13] mask_rev_in[14] mask_rev_in[15] mask_rev_in[16]
+ mask_rev_in[17] mask_rev_in[18] mask_rev_in[19] mask_rev_in[20]
+ mask_rev_in[21] mask_rev_in[22] mask_rev_in[23] mask_rev_in[24]
+ mask_rev_in[25] mask_rev_in[26] mask_rev_in[27] mask_rev_in[28]
+ mask_rev_in[29] mask_rev_in[30] mask_rev_in[31] pwr_ctrl_out[0]
+ pwr_ctrl_out[1] sram_ro_csb sram_ro_addr[0] reset serial_clock porb wb_rstn_i
+ sram_ro_addr[1] serial_resetn pwr_ctrl_out[3] pad_flash_clk VPWR pll_ena
+ pwr_ctrl_out[2] serial_load sram_ro_addr[2] sram_ro_addr[3] sram_ro_addr[4]
+ serial_data_1 sram_ro_addr[5] sram_ro_addr[6] serial_data_2 sram_ro_addr[7]
+ mgmt_gpio_in[0] sram_ro_clk sram_ro_data[0] mgmt_gpio_oeb[0] sram_ro_data[1]
+ sram_ro_data[2] mgmt_gpio_out[0] sram_ro_data[3] mgmt_gpio_in[1]
+ sram_ro_data[4] mgmt_gpio_in[4] sram_ro_data[5] mgmt_gpio_oeb[1]
+ sram_ro_data[6] sram_ro_data[7] mgmt_gpio_out[1] sram_ro_data[8]
+ mgmt_gpio_in[2] sram_ro_data[9] sram_ro_data[10] mgmt_gpio_oeb[2]
+ sram_ro_data[11] mgmt_gpio_out[2] sram_ro_data[12] mgmt_gpio_in[3]
+ sram_ro_data[13] sram_ro_data[14] sram_ro_data[15] mgmt_gpio_oeb[3]
+ sram_ro_data[16] mgmt_gpio_out[3] sram_ro_data[17] sram_ro_data[18]
+ sram_ro_data[19] sram_ro_data[20] mgmt_gpio_oeb[4] sram_ro_data[21]
+ mgmt_gpio_out[4] sram_ro_data[22] sram_ro_data[23] mgmt_gpio_in[5]
+ sram_ro_data[24] sram_ro_data[25] mgmt_gpio_oeb[5] sram_ro_data[26]
+ mgmt_gpio_out[5] sram_ro_data[27] sram_ro_data[28] mgmt_gpio_in[6]
+ sram_ro_data[29] sram_ro_data[30] mgmt_gpio_oeb[6] sram_ro_data[31]
+ mgmt_gpio_out[6] debug_in debug_mode mgmt_gpio_in[7] debug_oeb debug_out
+ mgmt_gpio_oeb[7] trap irq[0] mgmt_gpio_out[7] irq[1] mgmt_gpio_in[8] irq[2]
+ spi_sdoenb mgmt_gpio_oeb[8] spi_sdo mgmt_gpio_out[8] spi_sck wb_clk_i spi_csb
+ mgmt_gpio_in[9] spi_sdi ser_tx mgmt_gpio_oeb[9] ser_rx mgmt_gpio_out[9]
+ qspi_enabled uart_enabled mgmt_gpio_in[10] spi_enabled wb_ack_o
+ mgmt_gpio_oeb[10] wb_stb_i wb_dat_o[0] mgmt_gpio_out[10] wb_dat_o[1]
+ mgmt_gpio_in[11] wb_dat_o[2] wb_dat_o[3] mgmt_gpio_oeb[11] wb_dat_o[4]
+ mgmt_gpio_out[11] wb_dat_o[5] wb_dat_o[6] mgmt_gpio_in[12] wb_dat_o[7]
+ wb_dat_o[8] mgmt_gpio_oeb[12] wb_dat_o[9] mgmt_gpio_out[12] wb_dat_o[10]
+ wb_dat_o[11] mgmt_gpio_in[13] wb_dat_o[12] wb_dat_o[13] mgmt_gpio_oeb[13]
+ wb_dat_o[14] wb_dat_o[15] mgmt_gpio_out[13] wb_dat_o[16] mgmt_gpio_in[14]
+ wb_dat_o[17] wb_dat_o[18] mgmt_gpio_oeb[14] wb_dat_o[19] mgmt_gpio_out[14]
+ wb_dat_o[20] wb_dat_o[21] mgmt_gpio_in[15] wb_dat_o[22] wb_dat_o[23]
+ mgmt_gpio_oeb[15] wb_dat_o[24] mgmt_gpio_out[15] wb_dat_o[25] user_clock
+ wb_dat_o[26] mgmt_gpio_in[16] wb_dat_o[27] wb_dat_o[28] mgmt_gpio_oeb[16]
+ wb_dat_o[29] mgmt_gpio_out[33] mgmt_gpio_out[16] wb_dat_o[30] wb_dat_o[31]
+ mgmt_gpio_in[17] spimemio_flash_clk spimemio_flash_csb mgmt_gpio_out[17]
+ mgmt_gpio_oeb[17] spimemio_flash_io0_di spimemio_flash_io0_do
+ spimemio_flash_io0_oeb mgmt_gpio_out[32] mgmt_gpio_out[18] mgmt_gpio_in[18]
+ spimemio_flash_io1_di mgmt_gpio_out[31] mgmt_gpio_oeb[18]
+ spimemio_flash_io1_do mgmt_gpio_out[28] spimemio_flash_io1_oeb
+ spimemio_flash_io2_di mgmt_gpio_out[26] mgmt_gpio_out[30]
+ spimemio_flash_io2_do mgmt_gpio_out[20] mgmt_gpio_out[23] mgmt_gpio_in[19]
+ mgmt_gpio_out[19] mgmt_gpio_out[25] mgmt_gpio_out[37] wb_adr_i[3]
+ mgmt_gpio_out[21] mgmt_gpio_out[24] mgmt_gpio_out[27] mgmt_gpio_out[36]
+ mgmt_gpio_out[22] mgmt_gpio_out[29] spimemio_flash_io2_oeb
+ spimemio_flash_io3_do wb_adr_i[9] mgmt_gpio_out[34] wb_adr_i[0] wb_adr_i[6]
+ wb_we_i wb_adr_i[1] wb_adr_i[2] wb_adr_i[4] mgmt_gpio_in[37] wb_sel_i[3]
+ mgmt_gpio_oeb[28] mgmt_gpio_out[35] mgmt_gpio_oeb[37] mgmt_gpio_oeb[34]
+ mgmt_gpio_oeb[31] mgmt_gpio_oeb[36] spimemio_flash_io3_di mgmt_gpio_in[31]
+ spimemio_flash_io3_oeb wb_adr_i[8] wb_dat_i[10] wb_adr_i[5] wb_adr_i[7]
+ wb_adr_i[10] wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14] wb_adr_i[15]
+ wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19] wb_adr_i[20] wb_adr_i[21]
+ wb_adr_i[22] wb_adr_i[23] wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27]
+ wb_adr_i[28] wb_adr_i[29] wb_adr_i[30] wb_adr_i[31] wb_dat_i[0] wb_dat_i[1]
+ wb_dat_i[2] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6] wb_dat_i[7]
+ wb_dat_i[8] wb_dat_i[9] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13] wb_dat_i[14]
+ wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[20]
+ wb_dat_i[21] wb_dat_i[22] wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26]
+ wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[30] wb_dat_i[31] wb_sel_i[0]
+ wb_sel_i[1] wb_sel_i[2] wb_cyc_i usr1_vcc_pwrgood usr2_vcc_pwrgood
+ usr1_vdd_pwrgood usr2_vdd_pwrgood mgmt_gpio_in[20] mgmt_gpio_in[21]
+ mgmt_gpio_in[22] mgmt_gpio_in[23] mgmt_gpio_in[24] mgmt_gpio_in[25]
+ mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28] mgmt_gpio_in[29]
+ mgmt_gpio_in[30] mgmt_gpio_in[32] mgmt_gpio_in[33] mgmt_gpio_in[34]
+ mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_oeb[20] mgmt_gpio_oeb[21]
+ mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25]
+ mgmt_gpio_oeb[26] mgmt_gpio_oeb[27] mgmt_gpio_oeb[29] mgmt_gpio_oeb[30]
+ mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[35] mgmt_gpio_oeb[19] VGND
X$1 VPWR VGND pad_flash_clk_oeb VPWR \$96 VGND sky130_fd_sc_hd__buf_2
X$2 VPWR VGND pad_flash_csb VPWR \$136 VGND sky130_fd_sc_hd__buf_2
X$3 VPWR VGND pad_flash_csb_oeb VPWR \$97 VGND sky130_fd_sc_hd__buf_2
X$4 VPWR \$155 VGND VPWR pad_flash_io0_di VGND sky130_fd_sc_hd__clkbuf_1
X$5 VPWR VGND pad_flash_io0_do VPWR \$98 VGND sky130_fd_sc_hd__buf_2
X$6 VPWR VGND pad_flash_io0_ieb VPWR \$99 VGND sky130_fd_sc_hd__buf_2
X$7 VPWR VGND pad_flash_io0_oeb VPWR \$100 VGND sky130_fd_sc_hd__buf_2
X$8 VPWR VGND \$573 VPWR pad_flash_io1_di VGND sky130_fd_sc_hd__buf_2
X$9 VPWR VGND pad_flash_io1_do VPWR \$101 VGND sky130_fd_sc_hd__buf_2
X$10 VPWR VGND pad_flash_io1_ieb VPWR \$102 VGND sky130_fd_sc_hd__buf_2
X$11 VPWR VGND pad_flash_io1_oeb VPWR \$228 VGND sky130_fd_sc_hd__buf_2
X$12 VPWR VGND pll_dco_ena VPWR \$104 VGND sky130_fd_sc_hd__buf_2
X$13 VPWR VGND pll_div[0] VPWR \$105 VGND sky130_fd_sc_hd__buf_2
X$14 VPWR VGND pll_div[1] VPWR \$106 VGND sky130_fd_sc_hd__buf_2
X$15 VPWR VGND pll_div[2] VPWR \$107 VGND sky130_fd_sc_hd__buf_2
X$16 VPWR VGND pll_div[3] VPWR \$108 VGND sky130_fd_sc_hd__buf_2
X$17 VPWR VGND pll_div[4] VPWR \$109 VGND sky130_fd_sc_hd__buf_2
X$18 VPWR VGND pll_sel[0] VPWR \$137 VGND sky130_fd_sc_hd__buf_2
X$19 VPWR VGND pll_sel[1] VPWR \$110 VGND sky130_fd_sc_hd__buf_2
X$20 VPWR VGND pll_sel[2] VPWR \$111 VGND sky130_fd_sc_hd__buf_2
X$21 VPWR VGND pll90_sel[0] VPWR \$112 VGND sky130_fd_sc_hd__buf_2
X$22 VPWR VGND pll90_sel[1] VPWR \$113 VGND sky130_fd_sc_hd__buf_2
X$23 VPWR VGND pll90_sel[2] VPWR \$138 VGND sky130_fd_sc_hd__buf_2
X$24 VPWR VGND pll_trim[0] VPWR \$114 VGND sky130_fd_sc_hd__buf_2
X$25 VPWR VGND pll_trim[1] VPWR \$115 VGND sky130_fd_sc_hd__buf_2
X$26 VPWR VGND pll_trim[2] VPWR \$398 VGND sky130_fd_sc_hd__buf_2
X$27 VPWR VGND pll_trim[3] VPWR \$116 VGND sky130_fd_sc_hd__buf_2
X$28 VPWR VGND pll_trim[4] VPWR \$139 VGND sky130_fd_sc_hd__buf_2
X$29 VPWR VGND pll_trim[5] VPWR \$117 VGND sky130_fd_sc_hd__buf_2
X$30 VPWR VGND pll_trim[6] VPWR \$430 VGND sky130_fd_sc_hd__buf_2
X$31 VPWR VGND pll_trim[7] VPWR \$346 VGND sky130_fd_sc_hd__buf_2
X$32 VPWR VGND pll_trim[8] VPWR \$118 VGND sky130_fd_sc_hd__buf_2
X$33 VPWR VGND pll_trim[9] VPWR \$140 VGND sky130_fd_sc_hd__buf_2
X$34 VPWR VGND pll_trim[10] VPWR \$141 VGND sky130_fd_sc_hd__buf_2
X$35 VPWR VGND pll_trim[11] VPWR \$142 VGND sky130_fd_sc_hd__buf_2
X$36 VPWR VGND pll_trim[12] VPWR \$143 VGND sky130_fd_sc_hd__buf_2
X$37 VPWR VGND pll_trim[13] VPWR \$119 VGND sky130_fd_sc_hd__buf_2
X$38 VPWR VGND pll_trim[14] VPWR \$120 VGND sky130_fd_sc_hd__buf_2
X$39 VPWR VGND pll_trim[15] VPWR \$121 VGND sky130_fd_sc_hd__buf_2
X$40 VPWR VGND pll_trim[16] VPWR \$122 VGND sky130_fd_sc_hd__buf_2
X$41 VPWR VGND pll_trim[17] VPWR \$144 VGND sky130_fd_sc_hd__buf_2
X$42 VPWR VGND pll_trim[18] VPWR \$123 VGND sky130_fd_sc_hd__buf_2
X$43 VPWR VGND pll_trim[19] VPWR \$124 VGND sky130_fd_sc_hd__buf_2
X$44 VPWR VGND pll_trim[20] VPWR \$125 VGND sky130_fd_sc_hd__buf_2
X$45 VPWR VGND pll_trim[21] VPWR \$126 VGND sky130_fd_sc_hd__buf_2
X$46 VPWR VGND pll_trim[22] VPWR \$127 VGND sky130_fd_sc_hd__buf_2
X$47 VPWR VGND pll_trim[23] VPWR \$128 VGND sky130_fd_sc_hd__buf_2
X$48 VPWR VGND pll_trim[24] VPWR \$129 VGND sky130_fd_sc_hd__buf_2
X$49 VPWR VGND pll_trim[25] VPWR \$130 VGND sky130_fd_sc_hd__buf_2
X$50 VPWR VGND pll_bypass VPWR \$145 VGND sky130_fd_sc_hd__buf_2
X$51 VPWR \$156 VGND VPWR mask_rev_in[0] VGND sky130_fd_sc_hd__clkbuf_1
X$52 VPWR \$157 VGND VPWR mask_rev_in[1] VGND sky130_fd_sc_hd__clkbuf_1
X$53 VPWR \$158 VGND VPWR mask_rev_in[2] VGND sky130_fd_sc_hd__clkbuf_1
X$54 VPWR \$159 VGND VPWR mask_rev_in[3] VGND sky130_fd_sc_hd__clkbuf_1
X$55 VPWR \$160 VGND VPWR mask_rev_in[4] VGND sky130_fd_sc_hd__clkbuf_1
X$56 VPWR \$161 VGND VPWR mask_rev_in[5] VGND sky130_fd_sc_hd__clkbuf_1
X$57 VPWR \$162 VGND VPWR mask_rev_in[6] VGND sky130_fd_sc_hd__clkbuf_1
X$58 VPWR \$163 VGND VPWR mask_rev_in[7] VGND sky130_fd_sc_hd__clkbuf_1
X$59 VPWR VGND \$149 VPWR mask_rev_in[8] VGND sky130_fd_sc_hd__buf_2
X$60 VPWR \$89 VGND VPWR mask_rev_in[9] VGND sky130_fd_sc_hd__clkbuf_1
X$61 VPWR \$150 VGND VPWR mask_rev_in[10] VGND sky130_fd_sc_hd__clkbuf_1
X$62 VPWR \$164 VGND VPWR mask_rev_in[11] VGND sky130_fd_sc_hd__clkbuf_1
X$63 VPWR \$165 VGND VPWR mask_rev_in[12] VGND sky130_fd_sc_hd__clkbuf_1
X$64 VPWR \$94 VGND VPWR mask_rev_in[13] VGND sky130_fd_sc_hd__clkbuf_1
X$65 VPWR \$151 VGND VPWR mask_rev_in[14] VGND sky130_fd_sc_hd__clkbuf_1
X$66 VPWR \$146 VGND VPWR mask_rev_in[15] VGND sky130_fd_sc_hd__clkbuf_1
X$67 VPWR \$166 VGND VPWR mask_rev_in[16] VGND sky130_fd_sc_hd__clkbuf_1
X$68 VPWR \$167 VGND VPWR mask_rev_in[17] VGND sky130_fd_sc_hd__clkbuf_1
X$69 VPWR \$95 VGND VPWR mask_rev_in[18] VGND sky130_fd_sc_hd__clkbuf_1
X$70 VPWR \$168 VGND VPWR mask_rev_in[19] VGND sky130_fd_sc_hd__clkbuf_1
X$71 VPWR \$169 VGND VPWR mask_rev_in[20] VGND sky130_fd_sc_hd__clkbuf_1
X$72 VPWR \$170 VGND VPWR mask_rev_in[21] VGND sky130_fd_sc_hd__clkbuf_1
X$73 VPWR \$152 VGND VPWR mask_rev_in[22] VGND sky130_fd_sc_hd__clkbuf_1
X$74 VPWR \$171 VGND VPWR mask_rev_in[23] VGND sky130_fd_sc_hd__clkbuf_1
X$75 VPWR \$172 VGND VPWR mask_rev_in[24] VGND sky130_fd_sc_hd__clkbuf_1
X$76 VPWR \$173 VGND VPWR mask_rev_in[25] VGND sky130_fd_sc_hd__clkbuf_1
X$77 VPWR \$174 VGND VPWR mask_rev_in[26] VGND sky130_fd_sc_hd__clkbuf_1
X$78 VPWR \$175 VGND VPWR mask_rev_in[27] VGND sky130_fd_sc_hd__clkbuf_1
X$79 VPWR \$176 VGND VPWR mask_rev_in[28] VGND sky130_fd_sc_hd__clkbuf_1
X$80 VPWR \$153 VGND VPWR mask_rev_in[29] VGND sky130_fd_sc_hd__clkbuf_1
X$81 VPWR \$177 VGND VPWR mask_rev_in[30] VGND sky130_fd_sc_hd__clkbuf_1
X$82 VPWR \$178 VGND VPWR mask_rev_in[31] VGND sky130_fd_sc_hd__clkbuf_1
X$83 VPWR VGND pwr_ctrl_out[0] VPWR \$133 VGND sky130_fd_sc_hd__buf_2
X$84 VPWR VGND pwr_ctrl_out[1] VPWR \$134 VGND sky130_fd_sc_hd__buf_2
X$85 VPWR VGND sram_ro_csb VPWR \$91 VGND sky130_fd_sc_hd__buf_2
X$86 VPWR VGND sram_ro_addr[0] VPWR \$193 VGND sky130_fd_sc_hd__buf_2
X$87 VPWR VGND reset VPWR \$103 VGND sky130_fd_sc_hd__buf_2
X$88 VPWR VGND VPWR \$262 \$89 VGND sky130_fd_sc_hd__inv_2
X$89 VPWR serial_clock VGND VPWR \$147 VGND sky130_fd_sc_hd__clkbuf_1
X$90 VGND \$655 \$91 \$237 \$483 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_2
X$91 VGND \$493 \$91 \$183 \$523 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$92 VPWR VGND VPWR \$1164 \$91 VGND sky130_fd_sc_hd__inv_2
X$93 VGND porb \$655 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$94 VGND \$93 \$1369 \$5034 \$5107 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$95 VGND \$93 \$1452 \$5034 \$5018 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$96 VGND \$93 \$5079 \$5034 \$5378 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$97 VGND \$93 \$5495 \$5034 \$5426 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$98 VGND \$93 \$5423 \$5034 \$5416 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$99 VGND \$93 \$3831 \$5034 \$5338 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$100 VGND \$93 \$4897 \$5034 \$4921 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$101 VGND \$93 \$5432 \$5034 \$5431 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$102 VGND \$93 \$5215 \$5034 \$5407 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$103 VGND \$93 \$5681 \$5034 \$5693 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$104 VGND \$93 \$5686 \$5002 \$5669 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$105 VGND \$93 \$5610 \$5002 \$5716 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$106 VGND \$93 \$1550 \$1201 \$1832 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$107 VGND \$93 \$5116 \$5002 \$5176 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$108 VGND \$93 \$2070 \$1201 \$2092 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$109 VGND \$93 \$5176 \$5034 \$5306 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$110 VGND \$93 \$1324 \$1201 \$1674 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$111 VGND \$93 \$1398 \$1201 \$1935 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$112 VGND \$93 \$1636 \$1201 \$1635 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$113 VGND \$93 \$2244 \$1201 \$2260 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$114 VGND \$93 \$1488 \$1201 \$1849 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$115 VGND \$93 \$5531 \$5034 \$5545 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$116 VGND \$93 \$5748 \$5002 \$5763 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$117 VGND \$93 \$5651 \$5034 \$5670 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$118 VGND \$93 \$5648 \$5002 \$5761 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$119 VGND \$93 \$5204 \$5034 \$5163 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$120 VGND \$93 \$5226 \$5034 \$5260 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$121 VGND \$93 \$5649 \$5002 \$5700 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$122 VPWR VGND VPWR \$5235 \$93 VGND sky130_fd_sc_hd__inv_2
X$123 VGND \$93 \$5301 \$5034 \$5248 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$124 VGND wb_rstn_i \$93 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$125 VPWR VGND VPWR \$245 \$94 VGND sky130_fd_sc_hd__inv_2
X$126 VPWR VGND VPWR \$249 \$95 VGND sky130_fd_sc_hd__inv_2
X$127 VPWR \$96 VGND \$655 VPWR \$308 VGND sky130_fd_sc_hd__nor2_1
X$128 VPWR \$97 VGND \$655 VPWR \$235 VGND sky130_fd_sc_hd__nor2_1
X$129 VGND \$98 \$1395 \$780 \$235 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$130 VPWR VGND VPWR \$100 \$99 VGND sky130_fd_sc_hd__inv_2
X$131 VPWR \$99 VGND VPWR \$236 VGND sky130_fd_sc_hd__clkbuf_1
X$132 VPWR \$101 VGND VPWR \$225 VGND sky130_fd_sc_hd__clkbuf_1
X$133 VPWR VGND VPWR \$102 \$228 VGND sky130_fd_sc_hd__inv_2
X$134 VPWR VGND VPWR \$1654 \$103 VGND sky130_fd_sc_hd__inv_2
X$135 VPWR VGND \$103 VPWR \$865 VGND sky130_fd_sc_hd__buf_2
X$136 VGND \$280 \$104 \$293 \$273 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$137 VPWR VGND VPWR \$312 \$104 VGND sky130_fd_sc_hd__inv_2
X$138 VGND \$655 \$104 \$237 \$238 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$139 VPWR VGND VPWR \$389 \$105 VGND sky130_fd_sc_hd__inv_2
X$140 VPWR VGND \$202 \$183 \$105 \$212 \$195 VPWR VGND sky130_fd_sc_hd__a22o_1
X$141 VGND \$206 \$105 \$239 \$212 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$142 VGND \$655 \$106 \$239 \$332 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$143 VPWR VGND VPWR \$782 \$106 VGND sky130_fd_sc_hd__inv_2
X$144 VPWR VGND \$202 \$293 \$106 \$332 \$195 VPWR VGND sky130_fd_sc_hd__a22o_1
X$145 VPWR VGND VPWR \$360 \$107 VGND sky130_fd_sc_hd__inv_2
X$146 VGND \$206 \$107 \$239 \$313 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$147 VPWR VGND \$202 \$200 \$107 \$313 \$195 VPWR VGND sky130_fd_sc_hd__a22o_1
X$148 VPWR VGND VPWR \$314 \$108 VGND sky130_fd_sc_hd__inv_2
X$149 VPWR VGND \$202 \$281 \$108 \$240 \$195 VPWR VGND sky130_fd_sc_hd__a22o_1
X$150 VGND \$206 \$108 \$239 \$240 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$151 VGND \$206 \$109 \$239 \$203 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$152 VPWR \$274 \$109 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$153 VPWR VGND \$202 \$294 \$109 \$203 \$195 VPWR VGND sky130_fd_sc_hd__a22o_1
X$154 VPWR VGND VPWR \$557 \$110 VGND sky130_fd_sc_hd__inv_2
X$155 VGND \$655 \$110 \$239 \$538 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$156 VPWR VGND \$545 \$293 \$110 \$538 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$157 VGND \$655 \$111 \$239 \$683 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$158 VPWR VGND VPWR \$1017 \$111 VGND sky130_fd_sc_hd__inv_2
X$159 VPWR VGND \$545 \$200 \$111 \$683 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$160 VPWR VGND VPWR \$539 \$112 VGND sky130_fd_sc_hd__inv_2
X$161 VPWR VGND \$545 \$281 \$112 \$344 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$162 VGND \$206 \$112 \$241 \$344 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$163 VGND \$655 \$113 \$241 \$654 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_2
X$164 VPWR VGND VPWR \$1096 \$113 VGND sky130_fd_sc_hd__inv_2
X$165 VPWR VGND \$545 \$294 \$113 \$654 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$166 VPWR VGND VPWR \$333 \$114 VGND sky130_fd_sc_hd__inv_2
X$167 VGND \$206 \$114 \$241 \$220 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$168 VPWR VGND \$204 \$183 \$114 \$220 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$169 VPWR VGND VPWR \$334 \$115 VGND sky130_fd_sc_hd__inv_2
X$170 VGND \$206 \$115 \$241 \$275 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$171 VPWR VGND \$204 \$293 \$115 \$275 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$172 VPWR VGND VPWR \$335 \$116 VGND sky130_fd_sc_hd__inv_2
X$173 VGND \$206 \$116 \$241 \$270 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$174 VPWR VGND \$204 \$281 \$116 \$270 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$175 VPWR VGND \$204 \$184 \$117 \$213 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$176 VPWR VGND VPWR \$256 \$117 VGND sky130_fd_sc_hd__inv_2
X$177 VGND \$206 \$117 \$241 \$213 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$178 VPWR VGND VPWR \$412 \$118 VGND sky130_fd_sc_hd__inv_2
X$179 VGND \$206 \$118 \$196 \$362 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$180 VPWR VGND \$282 \$183 \$118 \$362 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$181 VPWR VGND VPWR \$284 \$119 VGND sky130_fd_sc_hd__inv_2
X$182 VGND \$206 \$119 \$196 \$242 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$183 VPWR VGND \$282 \$184 \$119 \$242 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$184 VPWR \$496 \$120 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$185 VGND \$206 \$120 \$196 \$447 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$186 VPWR VGND \$282 \$411 \$120 \$447 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$187 VPWR VGND VPWR \$185 \$121 VGND sky130_fd_sc_hd__inv_2
X$188 VGND \$206 \$121 \$196 \$317 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$189 VPWR VGND \$282 \$354 \$121 \$317 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$190 VPWR VGND VPWR \$364 \$122 VGND sky130_fd_sc_hd__inv_2
X$191 VGND \$206 \$122 \$198 \$199 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$192 VPWR VGND \$229 \$183 \$122 \$199 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$193 VPWR VGND VPWR \$214 \$123 VGND sky130_fd_sc_hd__inv_2
X$194 VGND \$206 \$123 \$198 \$186 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$195 VPWR VGND \$229 \$200 \$123 \$186 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$196 VPWR VGND VPWR \$295 \$124 VGND sky130_fd_sc_hd__inv_2
X$197 VGND \$206 \$124 \$198 \$231 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$198 VPWR VGND \$229 \$281 \$124 \$231 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$199 VPWR VGND VPWR \$476 \$125 VGND sky130_fd_sc_hd__inv_2
X$200 VGND \$206 \$125 \$198 \$404 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$201 VPWR VGND \$229 \$294 \$125 \$404 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$202 VPWR \$286 \$126 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$203 VGND \$206 \$126 \$198 \$257 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$204 VPWR VGND \$229 \$184 \$126 \$257 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$205 VPWR VGND VPWR \$403 \$127 VGND sky130_fd_sc_hd__inv_2
X$206 VGND \$206 \$127 \$198 \$383 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$207 VPWR VGND \$229 \$411 \$127 \$383 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$208 VPWR VGND VPWR \$498 \$128 VGND sky130_fd_sc_hd__inv_2
X$209 VGND \$206 \$128 \$198 \$425 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$210 VPWR VGND \$229 \$354 \$128 \$425 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$211 VGND \$208 \$129 \$183 \$277 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$212 VPWR VGND VPWR \$303 \$129 VGND sky130_fd_sc_hd__inv_2
X$213 VGND \$206 \$129 \$243 \$187 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$214 VGND \$357 \$130 \$293 \$277 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$215 VPWR VGND VPWR \$508 \$130 VGND sky130_fd_sc_hd__inv_2
X$216 VGND \$206 \$130 \$243 \$366 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$217 VGND \$132 \$254 \$453 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$218 VPWR VGND VPWR \$554 \$132 VGND sky130_fd_sc_hd__inv_2
X$219 VPWR VGND \$301 \$542 \$132 \$453 \$306 VPWR VGND sky130_fd_sc_hd__a22o_1
X$220 VPWR VGND pwr_ctrl_out[3] VPWR \$132 VGND sky130_fd_sc_hd__buf_2
X$221 VGND \$133 \$254 \$234 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$222 VPWR VGND \$133 \$269 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$223 VPWR VGND \$301 \$1171 \$133 \$234 \$306 VPWR VGND sky130_fd_sc_hd__a22o_1
X$224 VGND \$134 \$254 \$309 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$225 VPWR VGND VPWR \$1121 \$134 VGND sky130_fd_sc_hd__inv_2
X$226 VPWR VGND \$301 \$1179 \$134 \$309 \$306 VPWR VGND sky130_fd_sc_hd__a22o_1
X$227 VPWR VGND sram_ro_addr[1] VPWR \$182 VGND sky130_fd_sc_hd__buf_2
X$228 VGND \$136 \$1394 \$1333 \$235 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$229 VGND \$655 \$137 \$239 \$640 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$230 VPWR VGND VPWR \$1031 \$137 VGND sky130_fd_sc_hd__inv_2
X$231 VPWR VGND \$545 \$183 \$137 \$640 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$232 VPWR VGND VPWR \$615 \$138 VGND sky130_fd_sc_hd__inv_2
X$233 VPWR VGND \$545 \$184 \$138 \$558 \$525 VPWR VGND sky130_fd_sc_hd__a22o_1
X$234 VGND \$655 \$138 \$241 \$558 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$235 VPWR \$588 \$139 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$236 VGND \$206 \$139 \$241 \$474 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$237 VPWR VGND \$204 \$294 \$139 \$474 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$238 VGND \$206 \$140 \$196 \$197 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$239 VPWR VGND VPWR \$315 \$140 VGND sky130_fd_sc_hd__inv_2
X$240 VPWR VGND \$282 \$293 \$140 \$197 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$241 VPWR VGND VPWR \$507 \$141 VGND sky130_fd_sc_hd__inv_2
X$242 VGND \$206 \$141 \$196 \$446 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$243 VPWR VGND \$282 \$200 \$141 \$446 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$244 VPWR VGND VPWR \$316 \$142 VGND sky130_fd_sc_hd__inv_2
X$245 VGND \$206 \$142 \$196 \$276 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$246 VPWR VGND \$282 \$281 \$142 \$276 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$247 VPWR VGND VPWR \$338 \$143 VGND sky130_fd_sc_hd__inv_2
X$248 VPWR VGND \$282 \$294 \$143 \$207 \$283 VPWR VGND sky130_fd_sc_hd__a22o_1
X$249 VGND \$206 \$143 \$196 \$207 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$250 VPWR VGND VPWR \$527 \$144 VGND sky130_fd_sc_hd__inv_2
X$251 VGND \$206 \$144 \$196 \$378 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$252 VPWR VGND \$229 \$293 \$144 \$378 \$230 VPWR VGND sky130_fd_sc_hd__a22o_1
X$253 VGND \$946 \$145 \$183 \$1046 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$254 VPWR VGND VPWR \$1022 \$145 VGND sky130_fd_sc_hd__inv_2
X$255 VGND \$655 \$145 \$605 \$928 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$256 VPWR VGND VPWR \$263 \$146 VGND sky130_fd_sc_hd__inv_2
X$257 VPWR VGND \$745 VPWR \$695 \$147 VGND sky130_fd_sc_hd__nor2_2
X$258 VGND \$322 \$322 \$852 \$895 \$903 \$147 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_2
X$259 VPWR \$903 VPWR VGND \$1109 \$973 \$147 VGND sky130_fd_sc_hd__or3_2
X$260 VGND \$808 \$973 \$914 \$147 \$322 \$1011 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$261 VGND \$289 \$147 \$895 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$262 VGND \$147 \$534 \$694 \$300 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$263 VPWR VGND serial_resetn VPWR \$380 VGND sky130_fd_sc_hd__buf_2
X$264 VPWR \$1371 VPWR VGND \$1034 \$1329 \$149 VGND sky130_fd_sc_hd__or3b_1
X$265 VPWR VGND VPWR \$244 \$150 VGND sky130_fd_sc_hd__inv_2
X$266 VPWR VGND VPWR \$264 \$151 VGND sky130_fd_sc_hd__inv_2
X$267 VPWR VGND VPWR \$210 \$152 VGND sky130_fd_sc_hd__inv_2
X$268 VPWR \$255 \$153 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$269 VPWR \$328 VGND VPWR \$155 \$235 VGND sky130_fd_sc_hd__and2b_1
X$270 VPWR VGND VPWR \$258 \$156 VGND sky130_fd_sc_hd__inv_2
X$271 VPWR VGND VPWR \$285 \$157 VGND sky130_fd_sc_hd__inv_2
X$272 VPWR VGND \$158 \$488 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$273 VPWR VGND VPWR \$221 \$159 VGND sky130_fd_sc_hd__inv_2
X$274 VPWR VGND VPWR \$509 \$160 VGND sky130_fd_sc_hd__inv_2
X$275 VPWR VGND VPWR \$259 \$161 VGND sky130_fd_sc_hd__inv_2
X$276 VPWR VGND VPWR \$260 \$162 VGND sky130_fd_sc_hd__inv_2
X$277 VPWR VGND VPWR \$261 \$163 VGND sky130_fd_sc_hd__inv_2
X$278 VPWR VGND VPWR \$356 \$164 VGND sky130_fd_sc_hd__inv_2
X$279 VPWR VGND VPWR \$190 \$165 VGND sky130_fd_sc_hd__inv_2
X$280 VPWR VGND VPWR \$415 \$166 VGND sky130_fd_sc_hd__inv_2
X$281 VPWR VGND VPWR \$265 \$167 VGND sky130_fd_sc_hd__inv_2
X$282 VPWR \$215 \$168 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$283 VPWR VGND VPWR \$216 \$169 VGND sky130_fd_sc_hd__inv_2
X$284 VPWR \$217 \$170 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$285 VPWR VGND VPWR \$189 \$171 VGND sky130_fd_sc_hd__inv_2
X$286 VPWR VGND VPWR \$267 \$172 VGND sky130_fd_sc_hd__inv_2
X$287 VPWR \$253 \$173 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$288 VPWR \$763 \$174 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$289 VPWR \$563 \$175 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$290 VPWR \$635 \$176 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$291 VPWR VGND VPWR \$191 \$177 VGND sky130_fd_sc_hd__inv_2
X$292 VPWR \$764 \$178 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$293 VPWR pad_flash_clk VGND VPWR \$371 VGND sky130_fd_sc_hd__clkbuf_1
X$294 VPWR ser_tx VPWR VGND \$2620 VGND sky130_fd_sc_hd__buf_4
X$295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$297 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$298 VGND \$3483 \$3342 \$2996 \$1998 \$2336 \$3470 VPWR VPWR VGND
+ sky130_fd_sc_hd__a311oi_2
X$299 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$300 VPWR \$2336 \$3358 VGND \$3470 VPWR \$1962 VGND sky130_fd_sc_hd__nor3_1
X$301 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$302 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$303 VGND \$2410 \$3411 \$2678 \$4034 \$3248 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$306 VGND \$2929 \$3452 \$3471 \$3439 \$3100 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$307 VGND \$3153 \$3452 \$3440 \$3472 \$2817 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$308 VGND \$3154 \$3452 \$3440 \$3484 \$2680 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$310 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$311 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$312 VGND \$3259 \$3452 \$3485 \$3440 \$2874 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$313 VPWR \$3453 \$3259 VGND \$3432 VPWR \$3486 \$3473 VGND
+ sky130_fd_sc_hd__or4_2
X$314 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$315 VPWR \$3487 VGND \$3141 \$1963 VPWR VGND sky130_fd_sc_hd__or2_1
X$316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$317 VPWR \$3302 VGND \$3433 \$3474 VPWR VGND sky130_fd_sc_hd__or2_1
X$318 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$321 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$322 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$323 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$324 VPWR VGND \$3284 \$200 \$3475 \$3457 \$3304 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$331 VPWR VGND VPWR \$3435 \$3458 VGND sky130_fd_sc_hd__inv_2
X$332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$335 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$336 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$337 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$344 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$347 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$351 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$352 VPWR \$3488 VGND VPWR \$2247 \$2190 \$3476 \$2751 VGND
+ sky130_fd_sc_hd__o22a_1
X$353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$357 VGND \$3464 \$3526 \$3476 \$2544 \$2545 \$2400 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$358 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$359 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$360 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$361 VGND \$3477 \$3465 \$2497 \$1845 \$3478 \$1157 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$363 VPWR \$1423 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$364 VPWR \$3489 VGND VPWR \$1423 \$1966 \$3403 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$367 VPWR \$3479 VGND VPWR \$3168 \$2665 \$1601 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$368 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$371 VGND \$3466 \$3479 \$3480 \$2544 \$2545 \$3467 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$374 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$375 VPWR VGND VPWR \$3496 \$3408 VGND sky130_fd_sc_hd__inv_2
X$376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$377 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$380 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$382 VPWR VGND \$3169 \$411 \$3481 \$3490 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$383 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$384 VGND \$2989 \$3481 \$3425 \$3490 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$387 VPWR \$3482 VGND VPWR \$3468 VGND sky130_fd_sc_hd__clkbuf_1
X$388 VPWR VGND mgmt_gpio_oeb[9] VPWR \$3482 VGND sky130_fd_sc_hd__buf_2
X$389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$391 VPWR VGND ser_rx VPWR \$3094 VGND sky130_fd_sc_hd__buf_2
X$392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$394 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$396 VPWR \$2678 \$3499 \$2486 VPWR VGND \$3498 \$3255 VGND
+ sky130_fd_sc_hd__or4_1
X$397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$400 VGND \$3500 \$3341 \$3491 \$3099 \$3258 \$3501 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2111o_2
X$401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$402 VPWR VGND \$2873 \$3491 \$3502 VPWR \$3492 \$2941 VGND
+ sky130_fd_sc_hd__or4b_2
X$403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$405 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$406 VPWR \$3487 \$3504 VPWR \$3455 VGND VGND sky130_fd_sc_hd__and2_1
X$407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$408 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$409 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$410 VPWR \$3505 VGND \$3474 \$3362 VPWR VGND sky130_fd_sc_hd__or2_1
X$411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$412 VGND \$1850 \$3493 \$3506 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$413 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$415 VGND \$2777 \$3475 \$3413 \$3457 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$417 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$418 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$419 VPWR VGND VPWR \$3508 \$3475 VGND sky130_fd_sc_hd__inv_2
X$420 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$425 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$426 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$429 VGND \$3494 \$3522 \$1265 \$2525 \$2458 \$3537 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$431 VPWR \$3510 VGND VPWR \$1259 \$2724 \$3180 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$433 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$434 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$435 VGND \$3511 \$3494 \$2062 \$3495 \$3512 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$436 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$437 VGND \$3513 \$3509 \$2544 \$2545 \$2060 \$2063 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$438 VPWR \$3513 VGND VPWR \$3514 \$2665 \$3132 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$439 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$441 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$442 VPWR \$1730 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$443 VPWR \$3515 VGND VPWR \$1730 \$2665 \$3161 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$444 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$446 VGND \$3420 \$3515 \$3721 \$2544 \$2545 \$2841 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$449 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$451 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$452 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$456 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$457 VGND \$3901 \$3423 \$3496 \$2386 \$2614 \$3944 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$459 VGND \$3516 \$3489 \$3496 \$2043 \$1914 \$1880 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$460 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$463 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$464 VGND \$3424 \$3517 \$3518 \$2544 \$2545 \$2605 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$465 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$466 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$467 VPWR \$3477 VGND VPWR \$3519 \$1645 \$3467 \$2386 VGND
+ sky130_fd_sc_hd__o22a_1
X$468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$469 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$470 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$476 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$477 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$478 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$479 VPWR VGND \$3171 VPWR \$3520 VGND sky130_fd_sc_hd__clkbuf_4
X$480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$481 VPWR VGND \$3481 \$1856 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$485 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$486 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$489 VPWR spimemio_flash_csb VPWR VGND \$1394 VGND sky130_fd_sc_hd__buf_4
X$490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$492 VGND \$5145 \$5002 \$5492 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$493 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$495 VPWR \$4439 VPWR VGND \$5493 \$5482 VGND sky130_fd_sc_hd__or2_2
X$496 VGND \$4510 \$5493 \$5502 \$4833 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$497 VPWR \$5405 VPWR VGND \$4864 \$5502 \$5466 VGND sky130_fd_sc_hd__or3_1
X$498 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$499 VPWR \$5503 VGND \$5406 \$5147 VPWR VGND sky130_fd_sc_hd__or2_1
X$500 VPWR \$5509 VPWR VGND \$4833 \$4733 \$5406 VGND sky130_fd_sc_hd__or3_1
X$501 VGND \$5503 \$2571 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$502 VPWR \$5148 VGND \$5483 \$5494 VPWR VGND sky130_fd_sc_hd__or2_1
X$503 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$504 VGND \$4477 \$5469 \$5458 \$5471 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$506 VPWR \$5467 VGND \$5449 \$5246 VPWR \$5495 VGND sky130_fd_sc_hd__o21ai_2
X$507 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$508 VPWR \$5504 \$1078 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$511 VPWR \$5484 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$513 VPWR \$5511 VGND VPWR \$5484 VGND sky130_fd_sc_hd__clkbuf_1
X$514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$515 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$516 VPWR VGND \$5504 \$5496 \$5450 \$5441 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$518 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$520 VGND \$354 \$5486 \$1369 \$5531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$521 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$522 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$524 VGND \$2777 \$5473 \$5165 \$5472 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$526 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$527 VGND \$2777 \$5436 \$5165 \$5460 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$528 VPWR VGND \$5097 \$4774 \$5462 \$5451 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$530 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$531 VGND \$2777 \$5475 \$5408 \$5497 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$532 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$535 VPWR \$1077 \$5505 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$536 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$538 VPWR VGND \$5512 VPWR \$5239 VGND sky130_fd_sc_hd__clkbuf_4
X$539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$540 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$542 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$544 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$545 VPWR VGND \$5498 \$1171 \$5452 \$5476 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$546 VGND \$4761 \$5477 \$5367 \$5506 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$549 VPWR VGND \$5498 \$354 \$5499 \$5513 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$550 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$551 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$554 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$556 VGND \$3952 \$5272 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$557 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$558 VPWR VGND \$5500 \$3721 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$559 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$560 VGND \$4764 \$5479 \$5334 \$5489 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$561 VPWR VGND \$5344 \$1594 \$5480 \$5507 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$565 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$567 VPWR \$3247 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$568 VGND \$5515 \$3247 \$5501 \$3438 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$569 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$571 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$572 VGND \$5516 \$1594 \$5464 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$574 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$576 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$579 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$581 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$582 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$583 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$586 VPWR \$5404 VPWR VGND \$5517 \$5466 \$5519 VGND sky130_fd_sc_hd__or3b_1
X$587 VPWR \$5482 VGND \$5519 \$5517 VPWR VGND sky130_fd_sc_hd__or2_1
X$588 VPWR VGND VPWR \$5502 \$5517 VGND sky130_fd_sc_hd__inv_2
X$589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$590 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$592 VGND \$5509 \$5422 \$4833 \$5468 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$593 VPWR \$5468 VGND \$5406 \$4733 VPWR VGND sky130_fd_sc_hd__or2_1
X$594 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$595 VPWR VGND VPWR \$5469 \$5494 VGND sky130_fd_sc_hd__inv_2
X$596 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$597 VPWR \$5520 VPWR VGND \$5467 \$5471 \$5510 VGND sky130_fd_sc_hd__or3_2
X$598 VPWR \$5521 VPWR VGND \$5471 \$5510 \$5470 VGND sky130_fd_sc_hd__or3_1
X$599 VGND \$5521 \$4474 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$602 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$604 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$605 VGND \$5511 \$5496 \$4106 \$5522 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$608 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$609 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$612 VPWR \$4933 \$5523 VPWR \$3507 VGND VGND sky130_fd_sc_hd__and2_1
X$613 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$614 VPWR \$5533 VGND VPWR \$5523 VGND sky130_fd_sc_hd__clkbuf_1
X$615 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$616 VPWR VGND VPWR \$5270 \$5495 VGND sky130_fd_sc_hd__inv_2
X$617 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$618 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$619 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$620 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$622 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$626 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$627 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$629 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$630 VPWR VGND \$5388 \$1594 \$5475 \$5497 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$632 VGND \$2777 \$5505 \$5408 \$5524 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$635 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$636 VPWR VGND \$5546 \$3161 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$637 VPWR VGND \$5525 \$1594 \$5526 \$5535 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$638 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$639 VPWR VGND \$5526 \$2753 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$642 VPWR VGND \$5498 \$1594 \$5477 \$5506 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$644 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$647 VGND \$4761 \$5499 \$5367 \$5513 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$648 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$650 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$651 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$652 VPWR VGND \$5527 VPWR \$5264 VGND sky130_fd_sc_hd__clkbuf_4
X$653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$654 VGND \$4761 \$5488 \$5272 \$5487 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$655 VPWR VGND VPWR \$4558 \$5488 VGND sky130_fd_sc_hd__inv_2
X$656 VPWR VGND \$5344 \$1171 \$5500 \$5514 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$658 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$659 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$660 VGND \$4764 \$5480 \$5334 \$5507 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$662 VGND \$4764 \$5501 \$5334 \$5518 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$665 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$666 VPWR \$5549 VGND VPWR \$5516 \$4724 \$5528 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$668 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$669 VGND \$3952 \$5298 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$671 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$672 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$673 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$675 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$676 VPWR spi_sdoenb VPWR VGND \$3095 VGND sky130_fd_sc_hd__buf_4
X$677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$678 VPWR \$3094 VGND VPWR \$3080 VGND sky130_fd_sc_hd__clkbuf_1
X$679 VPWR \$3067 \$2857 \$3097 VPWR VGND \$3096 \$3068 VGND
+ sky130_fd_sc_hd__or4_1
X$680 VPWR VGND \$3057 VPWR \$3096 \$2320 VGND sky130_fd_sc_hd__nor2_2
X$681 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$682 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$683 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$685 VPWR \$3098 VGND \$2891 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$686 VPWR \$3099 VGND \$3098 \$3081 VPWR VGND sky130_fd_sc_hd__or2_1
X$687 VPWR \$3100 VGND \$3081 \$2352 VPWR VGND sky130_fd_sc_hd__or2_1
X$688 VPWR VGND VPWR \$3081 \$3069 VGND sky130_fd_sc_hd__inv_2
X$689 VGND \$2871 \$3069 \$3101 \$3082 \$2891 \$2700 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$690 VPWR \$3101 VGND \$2891 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$693 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$694 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$696 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$697 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$698 VPWR \$3102 VGND \$3083 \$2238 VPWR VGND sky130_fd_sc_hd__or2_1
X$699 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$701 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$702 VPWR VGND \$2775 \$200 \$3084 \$3103 \$2776 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$704 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$705 VGND \$856 \$3070 \$2556 \$3104 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$706 VPWR VGND \$2876 \$281 \$3070 \$3104 \$2934 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$707 VPWR VGND VPWR \$2876 \$2934 VGND sky130_fd_sc_hd__inv_2
X$708 VPWR VGND VPWR \$3071 \$3070 VGND sky130_fd_sc_hd__inv_2
X$709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$710 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$711 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$714 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$716 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$717 VPWR \$1570 VGND VPWR \$3106 \$1356 VGND sky130_fd_sc_hd__or2_4
X$718 VPWR \$3105 VGND VPWR \$2879 \$1954 \$2593 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$720 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$722 VGND \$3033 \$3120 \$684 \$785 \$2220 \$3071 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$727 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$728 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$729 VGND \$1868 \$3085 \$2908 \$2386 \$1340 \$3071 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$733 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$734 VGND \$1842 \$3147 \$3086 \$3087 VPWR \$2057 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$736 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$738 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$739 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$740 VPWR \$3108 VGND VPWR \$3089 \$1956 \$1915 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$743 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$744 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$745 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$746 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$747 VGND \$3109 \$3078 \$1823 \$2047 \$2048 \$3090 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$748 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$749 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$750 VGND \$3086 \$3091 \$3110 \$3149 \$1561 \$3092 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$753 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$754 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$755 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$756 VPWR \$3065 VGND VPWR \$3092 \$1966 \$3037 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$757 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$758 VPWR VGND VPWR \$3111 \$3049 VGND sky130_fd_sc_hd__inv_2
X$759 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$761 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$763 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$764 VPWR \$3112 \$3050 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$768 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$770 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$772 VPWR \$3066 VGND VPWR \$2829 VGND sky130_fd_sc_hd__clkbuf_1
X$773 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$774 VPWR VGND mgmt_gpio_oeb[8] VPWR \$3079 VGND sky130_fd_sc_hd__buf_2
X$775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$778 VPWR \$2551 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$779 VPWR \$1997 \$3080 VPWR \$2551 VGND VGND sky130_fd_sc_hd__and2_1
X$780 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$781 VPWR \$3139 VGND \$3068 \$3096 VPWR VGND sky130_fd_sc_hd__or2_1
X$782 VPWR \$3140 VGND \$3068 \$3098 VPWR VGND sky130_fd_sc_hd__or2_1
X$783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$784 VPWR \$3123 \$2892 \$3114 VPWR VGND \$3115 \$3098 VGND
+ sky130_fd_sc_hd__or4_1
X$785 VPWR \$3123 VGND \$2472 VPWR \$3124 VGND sky130_fd_sc_hd__nor2_1
X$786 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$788 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$789 VGND \$3082 \$3125 \$2741 \$3124 \$2700 \$3124 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$790 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$791 VPWR \$2741 \$3116 \$2514 \$2002 VGND \$2001 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$792 VPWR VPWR VGND \$3126 \$1376 VGND sky130_fd_sc_hd__clkbuf_2
X$793 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$795 VPWR \$3083 VGND \$2234 VPWR \$3155 VGND sky130_fd_sc_hd__nor2_1
X$796 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$797 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$798 VPWR \$3201 VGND \$3083 \$2259 VPWR VGND sky130_fd_sc_hd__or2_1
X$799 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$800 VPWR \$3142 VGND \$2258 VPWR \$3177 VGND sky130_fd_sc_hd__nor2_1
X$801 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$802 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$804 VGND \$2682 \$3117 \$2950 \$3083 \$3118 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$805 VPWR \$3119 VGND \$3118 \$2980 VPWR VGND sky130_fd_sc_hd__or2_1
X$806 VPWR \$3118 VGND \$2511 VPWR \$2949 VGND sky130_fd_sc_hd__nor2_1
X$807 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$808 VGND \$2777 \$3084 \$2556 \$3103 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$809 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$810 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$811 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$812 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$813 VPWR \$3127 VGND \$1340 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$814 VPWR VPWR VGND \$3127 \$2934 VGND sky130_fd_sc_hd__clkbuf_2
X$815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$817 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$818 VPWR VPWR VGND \$3128 \$2705 VGND sky130_fd_sc_hd__clkbuf_2
X$819 VPWR \$3128 VGND \$2384 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$820 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$821 VPWR \$1444 VGND VPWR \$3143 \$1342 VGND sky130_fd_sc_hd__or2_4
X$822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$823 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$824 VGND \$3120 \$3105 \$3129 \$2358 \$2274 \$3002 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$825 VGND \$3073 \$3130 \$1282 \$2525 \$2458 \$3131 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$828 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$829 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$832 VGND \$3145 \$2029 \$3144 \$1340 \$2384 \$3132 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$834 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$835 VPWR \$1570 VGND VPWR \$3121 \$1258 VGND sky130_fd_sc_hd__or2_4
X$836 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$837 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$838 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$843 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$844 VPWR \$3134 VGND VPWR \$2596 \$2559 \$2806 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$845 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$846 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$847 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$848 VPWR VPWR VGND \$3133 \$2808 VGND sky130_fd_sc_hd__clkbuf_2
X$849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$850 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$853 VGND \$3148 \$3135 \$3122 \$1715 \$1754 \$1023 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$854 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$855 VGND \$3110 \$1940 \$2906 \$1839 \$4239 \$3136 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$856 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$857 VPWR \$3209 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$858 VGND \$3091 \$2115 \$3137 \$3209 \$1879 \$1803 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$860 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$861 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$862 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$863 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$867 VPWR VGND \$2401 \$1171 \$3138 \$3151 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$870 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$872 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$874 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$875 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$876 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$877 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$878 VPWR VGND \$3213 \$2906 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$879 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$880 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$881 VPWR wb_adr_i[1] VPWR VGND \$4941 VGND sky130_fd_sc_hd__buf_4
X$882 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$883 VPWR VGND \$4916 VPWR wb_adr_i[0] VGND sky130_fd_sc_hd__clkbuf_4
X$884 VPWR wb_adr_i[2] VPWR VGND \$4942 VGND sky130_fd_sc_hd__buf_4
X$885 VPWR wb_adr_i[3] VPWR VGND \$5025 VGND sky130_fd_sc_hd__buf_4
X$886 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$887 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$888 VPWR wb_adr_i[4] VPWR VGND \$4881 VGND sky130_fd_sc_hd__buf_4
X$889 VPWR wb_adr_i[6] VPWR VGND \$4891 VGND sky130_fd_sc_hd__buf_4
X$890 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$891 VPWR \$5840 VPWR \$5841 \$5897 \$5813 \$5834 VGND VGND
+ sky130_fd_sc_hd__nand4_1
X$892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$893 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$894 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$895 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$896 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$897 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$898 VPWR \$5801 \$5883 VGND \$5884 VPWR \$5305 \$5770 VGND
+ sky130_fd_sc_hd__or4_2
X$899 VPWR \$5685 VGND \$5844 \$5845 VPWR VGND sky130_fd_sc_hd__or2_1
X$900 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$901 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$903 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$904 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$907 VGND \$5762 \$5917 \$5803 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$908 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$910 VGND \$5566 \$5918 \$5898 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$911 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$912 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$914 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$915 VPWR \$5423 \$5854 VPWR \$5908 VGND VGND sky130_fd_sc_hd__and2_1
X$916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$918 VGND \$5495 \$5079 \$5898 \$5909 \$5899 \$5900 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$920 VPWR \$5423 \$5909 VPWR \$5910 VGND VGND sky130_fd_sc_hd__and2_1
X$921 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$929 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$930 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$932 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$933 VGND \$5620 wb_sel_i[3] VPWR VPWR VGND sky130_fd_sc_hd__dlymetal6s2s_1
X$934 VPWR VPWR VGND wb_we_i \$5613 VGND sky130_fd_sc_hd__clkbuf_2
X$935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$936 VPWR VGND VPWR \$5911 \$1464 VGND sky130_fd_sc_hd__inv_4
X$937 VPWR VGND VPWR \$5912 \$1717 VGND sky130_fd_sc_hd__inv_4
X$938 VPWR \$4585 \$5913 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$939 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$940 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$941 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$943 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$944 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$945 VPWR \$5920 VGND VPWR \$5810 VGND sky130_fd_sc_hd__clkbuf_1
X$946 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$947 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$948 VPWR \$5921 VGND VPWR \$5811 VGND sky130_fd_sc_hd__clkbuf_1
X$949 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$950 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$952 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$953 VPWR \$5922 VGND VPWR \$5902 VGND sky130_fd_sc_hd__clkbuf_1
X$954 VPWR \$5902 VGND VPWR \$3037 VGND sky130_fd_sc_hd__clkbuf_1
X$955 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$956 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$957 VPWR \$5923 VGND VPWR \$5796 VGND sky130_fd_sc_hd__clkbuf_1
X$958 VGND \$5903 \$5932 \$4558 \$3636 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$959 VPWR VGND \$5914 \$3235 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$960 VPWR \$5924 VGND VPWR \$5890 VGND sky130_fd_sc_hd__clkbuf_1
X$961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$963 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$965 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$966 VPWR VGND mgmt_gpio_oeb[28] VPWR \$5831 VGND sky130_fd_sc_hd__buf_2
X$967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$968 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$969 VPWR \$5926 VGND VPWR \$1855 VGND sky130_fd_sc_hd__clkbuf_1
X$970 VPWR \$5927 VGND VPWR \$5926 VGND sky130_fd_sc_hd__clkbuf_1
X$971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$972 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$973 VPWR VGND VPWR \$4498 \$5915 VGND sky130_fd_sc_hd__inv_2
X$974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$975 VPWR \$5928 VGND VPWR \$5798 VGND sky130_fd_sc_hd__clkbuf_1
X$976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$977 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$978 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$979 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$980 VPWR \$5823 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$983 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$984 VPWR \$5904 VGND VPWR \$3092 VGND sky130_fd_sc_hd__clkbuf_1
X$985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$987 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$990 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$991 VPWR VGND mgmt_gpio_out[35] VPWR \$5412 VGND sky130_fd_sc_hd__buf_2
X$992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$993 VPWR VGND mgmt_gpio_oeb[37] VPWR \$5903 VGND sky130_fd_sc_hd__buf_2
X$994 VPWR mgmt_gpio_in[37] VPWR VGND \$5616 VGND sky130_fd_sc_hd__buf_4
X$995 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$996 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$998 VPWR \$5823 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$999 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1000 VPWR VGND \$5932 VPWR spimemio_flash_io3_oeb VGND sky130_fd_sc_hd__buf_2
X$1001 VGND wb_adr_i[5] \$4864 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1002 VPWR \$5872 VGND VPWR wb_adr_i[8] VGND sky130_fd_sc_hd__clkbuf_1
X$1003 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1004 VGND wb_adr_i[7] \$4853 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1005 VPWR VGND spimemio_flash_io3_di VPWR \$5882 VGND sky130_fd_sc_hd__buf_2
X$1006 VPWR \$5813 VGND VPWR wb_adr_i[10] VGND sky130_fd_sc_hd__clkbuf_1
X$1007 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1008 VPWR \$5841 VGND VPWR wb_adr_i[11] VGND sky130_fd_sc_hd__clkbuf_1
X$1009 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1010 VPWR \$5840 VGND VPWR wb_adr_i[12] VGND sky130_fd_sc_hd__clkbuf_1
X$1011 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1013 VPWR \$5834 VGND VPWR wb_adr_i[13] VGND sky130_fd_sc_hd__clkbuf_1
X$1014 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1015 VPWR \$5815 VGND VPWR wb_adr_i[14] VGND sky130_fd_sc_hd__clkbuf_1
X$1016 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1017 VPWR \$5842 VGND VPWR wb_adr_i[15] VGND sky130_fd_sc_hd__clkbuf_1
X$1018 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1019 VPWR \$5835 VGND VPWR wb_adr_i[16] VGND sky130_fd_sc_hd__clkbuf_1
X$1020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1021 VPWR \$5825 VGND VPWR wb_adr_i[17] VGND sky130_fd_sc_hd__clkbuf_1
X$1022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1023 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1024 VPWR \$5843 VGND VPWR wb_adr_i[18] VGND sky130_fd_sc_hd__clkbuf_1
X$1025 VPWR \$5875 VGND VPWR wb_adr_i[19] VGND sky130_fd_sc_hd__clkbuf_1
X$1026 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1027 VPWR VGND \$5684 VPWR wb_adr_i[20] VGND sky130_fd_sc_hd__buf_2
X$1028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1029 VPWR VGND \$5659 VPWR wb_adr_i[21] VGND sky130_fd_sc_hd__buf_2
X$1030 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1031 VPWR \$5844 VGND VPWR wb_adr_i[22] VGND sky130_fd_sc_hd__clkbuf_1
X$1032 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1033 VPWR \$5845 VGND VPWR wb_adr_i[23] VGND sky130_fd_sc_hd__clkbuf_1
X$1034 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1035 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1036 VPWR \$5846 VGND VPWR wb_adr_i[24] VGND sky130_fd_sc_hd__clkbuf_1
X$1037 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1038 VPWR \$5876 VGND VPWR wb_adr_i[25] VGND sky130_fd_sc_hd__clkbuf_1
X$1039 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1040 VPWR \$5847 VGND VPWR wb_adr_i[26] VGND sky130_fd_sc_hd__clkbuf_1
X$1041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1042 VPWR \$5849 VGND VPWR wb_adr_i[27] VGND sky130_fd_sc_hd__clkbuf_1
X$1043 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1044 VPWR \$5816 VGND VPWR wb_adr_i[28] VGND sky130_fd_sc_hd__clkbuf_1
X$1045 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1046 VPWR \$5848 VGND VPWR wb_adr_i[29] VGND sky130_fd_sc_hd__clkbuf_1
X$1047 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1049 VPWR \$5817 VGND VPWR wb_adr_i[30] VGND sky130_fd_sc_hd__clkbuf_1
X$1050 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1051 VPWR \$5850 VGND VPWR wb_adr_i[31] VGND sky130_fd_sc_hd__clkbuf_1
X$1052 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1053 VPWR \$5934 VGND VPWR wb_dat_i[0] VGND sky130_fd_sc_hd__clkbuf_1
X$1054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1055 VPWR \$5885 VGND VPWR wb_dat_i[1] VGND sky130_fd_sc_hd__clkbuf_1
X$1056 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1057 VPWR \$5917 VGND VPWR wb_dat_i[2] VGND sky130_fd_sc_hd__clkbuf_1
X$1058 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1059 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1060 VPWR \$5886 VGND VPWR wb_dat_i[3] VGND sky130_fd_sc_hd__clkbuf_1
X$1061 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1062 VPWR \$5791 VGND VPWR wb_dat_i[4] VGND sky130_fd_sc_hd__clkbuf_1
X$1063 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1064 VPWR \$5826 VGND VPWR wb_dat_i[5] VGND sky130_fd_sc_hd__clkbuf_1
X$1065 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1066 VPWR \$5792 VGND VPWR wb_dat_i[6] VGND sky130_fd_sc_hd__clkbuf_1
X$1067 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1068 VPWR \$5918 VGND VPWR wb_dat_i[7] VGND sky130_fd_sc_hd__clkbuf_1
X$1069 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1070 VPWR \$5852 VGND VPWR wb_dat_i[8] VGND sky130_fd_sc_hd__clkbuf_1
X$1071 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1072 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1073 VPWR \$5935 VGND VPWR wb_dat_i[9] VGND sky130_fd_sc_hd__clkbuf_1
X$1074 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1075 VPWR \$5782 VGND VPWR wb_dat_i[10] VGND sky130_fd_sc_hd__clkbuf_1
X$1076 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1077 VPWR \$5936 VGND VPWR wb_dat_i[11] VGND sky130_fd_sc_hd__clkbuf_1
X$1078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1079 VPWR \$5878 VGND VPWR wb_dat_i[12] VGND sky130_fd_sc_hd__clkbuf_1
X$1080 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1081 VPWR \$5785 VGND VPWR wb_dat_i[13] VGND sky130_fd_sc_hd__clkbuf_1
X$1082 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1083 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1084 VPWR \$5827 VGND VPWR wb_dat_i[14] VGND sky130_fd_sc_hd__clkbuf_1
X$1085 VPWR \$5899 VGND VPWR wb_dat_i[15] VGND sky130_fd_sc_hd__clkbuf_1
X$1086 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1087 VPWR \$5756 VGND VPWR wb_dat_i[16] VGND sky130_fd_sc_hd__clkbuf_1
X$1088 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1089 VPWR \$5908 VGND VPWR wb_dat_i[17] VGND sky130_fd_sc_hd__clkbuf_1
X$1090 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1091 VPWR \$5783 VGND VPWR wb_dat_i[18] VGND sky130_fd_sc_hd__clkbuf_1
X$1092 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1093 VPWR \$5860 VGND VPWR wb_dat_i[19] VGND sky130_fd_sc_hd__clkbuf_1
X$1094 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1095 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1096 VPWR \$5861 VGND VPWR wb_dat_i[20] VGND sky130_fd_sc_hd__clkbuf_1
X$1097 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1098 VPWR \$5862 VGND VPWR wb_dat_i[21] VGND sky130_fd_sc_hd__clkbuf_1
X$1099 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1100 VPWR \$5787 VGND VPWR wb_dat_i[22] VGND sky130_fd_sc_hd__clkbuf_1
X$1101 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1102 VPWR \$5910 VGND VPWR wb_dat_i[23] VGND sky130_fd_sc_hd__clkbuf_1
X$1103 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1104 VPWR \$5853 VGND VPWR wb_dat_i[24] VGND sky130_fd_sc_hd__clkbuf_1
X$1105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1106 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1107 VPWR \$5855 VGND VPWR wb_dat_i[25] VGND sky130_fd_sc_hd__clkbuf_1
X$1108 VPWR \$5765 VGND VPWR wb_dat_i[26] VGND sky130_fd_sc_hd__clkbuf_1
X$1109 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1110 VPWR \$5856 VGND VPWR wb_dat_i[27] VGND sky130_fd_sc_hd__clkbuf_1
X$1111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1112 VPWR \$5858 VGND VPWR wb_dat_i[28] VGND sky130_fd_sc_hd__clkbuf_1
X$1113 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1114 VPWR \$5786 VGND VPWR wb_dat_i[29] VGND sky130_fd_sc_hd__clkbuf_1
X$1115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1116 VPWR \$5859 VGND VPWR wb_dat_i[30] VGND sky130_fd_sc_hd__clkbuf_1
X$1117 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1118 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1119 VPWR \$5900 VGND VPWR wb_dat_i[31] VGND sky130_fd_sc_hd__clkbuf_1
X$1120 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1121 VPWR \$5701 VGND VPWR wb_sel_i[0] VGND sky130_fd_sc_hd__clkbuf_1
X$1122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1123 VPWR \$5688 VGND VPWR wb_sel_i[1] VGND sky130_fd_sc_hd__clkbuf_1
X$1124 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1125 VGND \$5614 wb_sel_i[2] VPWR VPWR VGND sky130_fd_sc_hd__dlymetal6s2s_1
X$1126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1129 VGND \$5837 wb_cyc_i VPWR VPWR VGND sky130_fd_sc_hd__dlymetal6s2s_1
X$1130 VPWR \$5913 VGND VPWR usr1_vcc_pwrgood VGND sky130_fd_sc_hd__clkbuf_1
X$1131 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1132 VPWR \$5788 VGND VPWR usr2_vcc_pwrgood VGND sky130_fd_sc_hd__clkbuf_1
X$1133 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1134 VPWR \$5912 VGND VPWR usr1_vdd_pwrgood VGND sky130_fd_sc_hd__clkbuf_1
X$1135 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1136 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1137 VPWR \$5911 VGND VPWR usr2_vdd_pwrgood VGND sky130_fd_sc_hd__clkbuf_1
X$1138 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1139 VPWR VPWR VGND mgmt_gpio_in[20] \$5702 VGND sky130_fd_sc_hd__clkbuf_2
X$1140 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1141 VPWR VGND mgmt_gpio_oeb[20] VPWR \$5888 VGND sky130_fd_sc_hd__buf_2
X$1142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1143 VPWR VGND \$3969 VPWR mgmt_gpio_in[21] VGND sky130_fd_sc_hd__clkbuf_4
X$1144 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1145 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1146 VPWR VGND mgmt_gpio_oeb[21] VPWR \$5889 VGND sky130_fd_sc_hd__buf_2
X$1147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1148 VPWR VGND \$4232 VPWR mgmt_gpio_in[22] VGND sky130_fd_sc_hd__clkbuf_4
X$1149 VPWR VGND mgmt_gpio_oeb[22] VPWR \$5920 VGND sky130_fd_sc_hd__buf_2
X$1150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1151 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1152 VPWR VPWR VGND mgmt_gpio_in[23] \$5134 VGND sky130_fd_sc_hd__clkbuf_2
X$1153 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1154 VPWR VGND mgmt_gpio_oeb[23] VPWR \$5921 VGND sky130_fd_sc_hd__buf_2
X$1155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1156 VPWR \$5863 VGND VPWR mgmt_gpio_in[24] VGND sky130_fd_sc_hd__clkbuf_1
X$1157 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1158 VPWR VGND mgmt_gpio_oeb[24] VPWR \$5922 VGND sky130_fd_sc_hd__buf_2
X$1159 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1160 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1161 VPWR VGND \$3948 VPWR mgmt_gpio_in[25] VGND sky130_fd_sc_hd__clkbuf_4
X$1162 VPWR VGND mgmt_gpio_oeb[25] VPWR \$5923 VGND sky130_fd_sc_hd__buf_2
X$1163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1164 VPWR \$5914 VGND VPWR mgmt_gpio_in[26] VGND sky130_fd_sc_hd__clkbuf_1
X$1165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1166 VPWR VGND mgmt_gpio_oeb[26] VPWR \$5924 VGND sky130_fd_sc_hd__buf_2
X$1167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1168 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1169 VPWR \$5865 VGND VPWR mgmt_gpio_in[27] VGND sky130_fd_sc_hd__clkbuf_1
X$1170 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1171 VPWR VGND mgmt_gpio_oeb[27] VPWR \$5797 VGND sky130_fd_sc_hd__buf_2
X$1172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1173 VGND \$5940 mgmt_gpio_in[28] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$1174 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1175 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1176 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1177 VGND \$5941 mgmt_gpio_in[29] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$1178 VPWR VGND mgmt_gpio_oeb[29] VPWR \$5927 VGND sky130_fd_sc_hd__buf_2
X$1179 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1180 VPWR \$5915 VGND VPWR mgmt_gpio_in[30] VGND sky130_fd_sc_hd__clkbuf_1
X$1181 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1182 VPWR VGND mgmt_gpio_oeb[30] VPWR \$5928 VGND sky130_fd_sc_hd__buf_2
X$1183 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1184 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1185 VGND \$5929 \$5823 \$5722 \$3636 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1186 VPWR VGND mgmt_gpio_oeb[31] VPWR \$5891 VGND sky130_fd_sc_hd__buf_2
X$1187 VPWR \$5866 VGND VPWR mgmt_gpio_in[31] VGND sky130_fd_sc_hd__clkbuf_1
X$1188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1189 VPWR VGND \$3588 VPWR mgmt_gpio_in[32] VGND sky130_fd_sc_hd__clkbuf_4
X$1190 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1191 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1192 VPWR VGND mgmt_gpio_oeb[32] VPWR \$5892 VGND sky130_fd_sc_hd__buf_2
X$1193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1194 VPWR VGND \$3755 VPWR mgmt_gpio_in[33] VGND sky130_fd_sc_hd__clkbuf_4
X$1195 VPWR VGND mgmt_gpio_oeb[33] VPWR \$5893 VGND sky130_fd_sc_hd__buf_2
X$1196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1197 VPWR VGND mgmt_gpio_oeb[34] VPWR \$5812 VGND sky130_fd_sc_hd__buf_2
X$1198 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1199 VGND mgmt_gpio_in[34] \$3429 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1200 VPWR \$5867 VGND VPWR mgmt_gpio_in[35] VGND sky130_fd_sc_hd__clkbuf_1
X$1201 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1202 VPWR VGND mgmt_gpio_oeb[35] VPWR \$4926 VGND sky130_fd_sc_hd__buf_2
X$1203 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1204 VPWR VGND mgmt_gpio_oeb[36] VPWR \$5887 VGND sky130_fd_sc_hd__buf_2
X$1205 VPWR VGND mgmt_gpio_oeb[19] VPWR \$5894 VGND sky130_fd_sc_hd__buf_2
X$1206 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1207 VPWR mgmt_gpio_in[36] VPWR VGND \$5595 VGND sky130_fd_sc_hd__buf_4
X$1208 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1210 VGND spimemio_flash_io1_do \$225 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1212 VPWR \$5667 VGND VPWR \$5358 \$5439 \$5448 \$1769 VGND
+ sky130_fd_sc_hd__o22a_1
X$1213 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1214 VPWR \$5668 VGND VPWR \$5403 \$5439 \$1619 \$5448 VGND
+ sky130_fd_sc_hd__o22a_1
X$1215 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1217 VPWR \$5647 VGND \$5632 \$5466 VPWR \$5646 VGND sky130_fd_sc_hd__o21ai_2
X$1218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1220 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1221 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1222 VGND \$5659 \$5618 \$5483 \$5471 \$5683 \$5678 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$1223 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1224 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1226 VGND \$5660 \$2015 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$1227 VPWR \$5661 VPWR VGND \$4603 VGND sky130_fd_sc_hd__buf_4
X$1228 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1230 VPWR \$5669 VGND VPWR \$5662 VGND sky130_fd_sc_hd__clkbuf_1
X$1231 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1232 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1233 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1234 VGND \$3732 \$5450 \$1369 \$5748 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$1235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1236 VPWR \$5670 VGND VPWR \$5680 VGND sky130_fd_sc_hd__clkbuf_1
X$1237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1238 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1239 VGND \$4023 \$780 \$1369 \$5681 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$1240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1241 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1242 VPWR VGND \$5192 \$3694 \$5663 \$5671 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1246 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1249 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1251 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1252 VPWR VGND \$5388 \$411 \$5656 \$5672 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1253 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1254 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1255 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1256 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1257 VPWR \$4670 \$5656 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1259 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1261 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1262 VPWR VGND \$5525 \$411 \$5629 \$5673 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1263 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1264 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1265 VGND \$2777 \$5629 \$5367 \$5673 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1269 VPWR VGND \$5498 \$184 \$5657 \$5674 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1270 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1272 VPWR VGND \$5657 \$3478 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$1273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1277 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1280 VPWR VGND \$5627 \$1594 \$5664 \$5644 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1281 VGND \$5664 \$1373 mgmt_gpio_out[28] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$1282 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1285 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1287 VPWR VGND \$5345 \$1594 \$5658 \$5645 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1289 VGND \$4764 \$5652 \$5298 \$5650 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$1290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1291 VPWR VGND \$5335 \$184 \$5665 \$5676 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1293 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1294 VPWR VGND \$5335 \$3694 \$5666 \$5677 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1297 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1298 VPWR VGND mgmt_gpio_oeb[18] VPWR \$5653 VGND sky130_fd_sc_hd__buf_2
X$1299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1301 VGND \$5358 \$5002 \$5667 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$1302 VGND \$5403 \$5002 \$5668 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$1303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1306 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1309 VPWR VGND VPWR \$5690 \$5682 VGND sky130_fd_sc_hd__inv_2
X$1310 VPWR VGND VPWR \$5678 \$5683 VGND sky130_fd_sc_hd__inv_2
X$1311 VPWR \$5494 VGND VPWR \$5684 \$5683 \$5679 \$5678 VGND
+ sky130_fd_sc_hd__o22a_1
X$1312 VPWR VGND \$5690 \$5618 \$5659 \$5510 \$5682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1313 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1314 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1315 VPWR \$5661 VPWR VGND \$5659 \$5679 \$5685 VGND sky130_fd_sc_hd__or3_1
X$1316 VPWR \$5660 VPWR VGND \$5659 \$5684 \$5685 VGND sky130_fd_sc_hd__or3_1
X$1317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1318 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1319 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1321 VGND \$5662 \$5686 \$5691 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1322 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1323 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1324 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1326 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1327 VGND \$5680 \$5651 \$5692 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1328 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1329 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1330 VPWR \$5558 VGND VPWR \$5687 VGND sky130_fd_sc_hd__clkbuf_1
X$1331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1332 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1333 VPWR \$5613 \$5586 VPWR \$5688 VGND VGND sky130_fd_sc_hd__and2_1
X$1334 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1335 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1336 VGND \$2777 \$5663 \$5165 \$5671 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$1337 VGND \$5663 \$1925 VPWR VPWR VGND sky130_fd_sc_hd__inv_8
X$1338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1339 VPWR VGND \$5689 \$2896 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$1340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1341 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1342 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1344 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1345 VGND \$2777 \$5656 \$5408 \$5672 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1348 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1349 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1351 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1355 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1356 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1358 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1359 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1360 VGND \$4761 \$5657 \$5367 \$5674 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1363 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1365 VGND \$5630 \$1320 mgmt_gpio_out[25] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$1366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1367 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1369 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1370 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1372 VGND \$4764 \$5698 \$5334 \$5694 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1376 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1377 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1378 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1380 VGND \$4764 \$5665 \$5298 \$5676 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1381 VGND \$4764 \$5666 \$5298 \$5677 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1382 VGND \$5695 \$3694 \$5666 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1383 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1384 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1386 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1387 VGND spi_sdo \$3172 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1391 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1392 VPWR \$3198 VGND \$3067 \$3123 VPWR VGND sky130_fd_sc_hd__or2_1
X$1393 VPWR \$3115 VGND \$3124 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$1394 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1395 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1396 VPWR VGND VPWR \$3173 \$3101 VGND sky130_fd_sc_hd__inv_2
X$1397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1399 VPWR \$2741 \$3174 \$2659 \$1999 VGND \$2001 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$1400 VPWR \$1919 \$3199 \$2795 VPWR VGND \$3174 \$3153 VGND
+ sky130_fd_sc_hd__or4_1
X$1401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1402 VPWR \$2041 \$3175 \$2714 VPWR VGND \$3116 \$3154 VGND
+ sky130_fd_sc_hd__or4_1
X$1403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1404 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1406 VPWR \$3156 VGND \$2336 \$3155 VPWR VGND sky130_fd_sc_hd__or2_1
X$1407 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1408 VPWR VPWR VGND \$3156 \$3141 VGND sky130_fd_sc_hd__clkbuf_2
X$1409 VGND \$2223 \$3157 \$3201 \$3176 \$3177 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$1410 VPWR VPWR \$2996 VGND \$3141 \$3178 \$3142 VGND sky130_fd_sc_hd__o21ai_1
X$1411 VPWR \$3177 VGND \$3141 VPWR \$1897 VGND sky130_fd_sc_hd__nor2_1
X$1412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1413 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1414 VPWR \$3179 VGND \$3176 \$3102 VPWR VGND sky130_fd_sc_hd__or2_1
X$1415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1417 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1418 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1420 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1421 VPWR \$3180 \$3084 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1424 VPWR VGND \$2876 \$200 \$3158 \$3202 \$2934 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1426 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1427 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1429 VPWR VGND \$2703 \$200 \$3159 \$3215 \$2705 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1430 VPWR VGND VPWR \$2703 \$2705 VGND sky130_fd_sc_hd__inv_2
X$1431 VPWR \$1570 VGND VPWR \$3181 \$1444 VGND sky130_fd_sc_hd__or2_4
X$1432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1433 VPWR VGND VPWR \$3183 \$2869 VGND sky130_fd_sc_hd__inv_2
X$1434 VGND \$3203 \$3182 \$3307 \$3143 \$686 \$812 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1435 VGND \$3184 \$1034 \$1258 \$3183 \$3143 \$3563 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$1436 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1437 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1438 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1439 VPWR \$3130 VGND VPWR \$3071 \$2456 \$2999 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$1440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1442 VGND \$3034 \$3160 \$3035 \$2116 \$1536 \$1817 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1444 VPWR \$1588 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1445 VGND \$3182 \$1763 \$3107 \$1588 \$1034 \$1356 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1447 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1448 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1449 VGND \$2787 \$3184 \$2936 \$2314 \$1625 \$3161 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1450 VGND \$3205 \$1865 \$819 \$1507 \$3121 \$3162 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1451 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1452 VGND \$3164 \$3163 \$2863 \$2751 \$2366 \$2983 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1454 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1455 VPWR VGND VPWR \$3147 \$3146 \$3165 \$3185 \$3164 VGND
+ sky130_fd_sc_hd__and4_1
X$1456 VGND \$3206 \$3166 \$3235 \$4239 \$1114 \$747 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1457 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1458 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1459 VPWR \$3166 VGND VPWR \$646 \$1507 \$2449 \$1867 VGND
+ sky130_fd_sc_hd__o22a_1
X$1460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1461 VGND \$3208 \$3134 \$2666 \$2750 \$2541 \$2587 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1463 VGND \$3187 \$3186 \$758 \$1953 \$1987 \$3089 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1464 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1465 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1466 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1467 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1468 VGND \$3189 \$1560 \$1847 \$3167 \$2375 \$3188 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$1469 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1471 VPWR \$3135 VGND VPWR \$1320 \$1776 \$1925 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$1472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1474 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1475 VPWR \$3191 VGND VPWR \$3111 \$2325 \$3168 \$1676 VGND
+ sky130_fd_sc_hd__o22a_1
X$1476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1477 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1478 VPWR \$3190 VGND VPWR \$620 \$2045 \$3038 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$1479 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1480 VGND \$3193 \$3466 \$3192 \$3048 VPWR \$983 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$1481 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1482 VPWR VGND VPWR \$3194 \$1997 VGND sky130_fd_sc_hd__inv_2
X$1483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1484 VPWR VGND \$2401 \$354 \$3150 \$3229 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1486 VPWR \$3195 VGND \$1879 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$1487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1488 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1489 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1490 VGND \$2989 \$3138 \$2450 \$3151 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$1491 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1492 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1493 VPWR VGND VPWR \$2502 \$3170 VGND sky130_fd_sc_hd__inv_2
X$1494 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1495 VPWR VGND \$3169 \$1594 \$3170 \$3196 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1497 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1500 VGND \$1152 \$3213 \$2232 \$3197 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1502 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1503 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1505 VPWR \$3340 \$2656 \$3332 VPWR VGND \$3198 \$3140 VGND
+ sky130_fd_sc_hd__or4_1
X$1506 VPWR \$3231 VPWR VGND \$3115 \$3096 \$3198 VGND sky130_fd_sc_hd__or3_1
X$1507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1511 VPWR VGND \$2002 VPWR \$3230 VGND sky130_fd_sc_hd__buf_2
X$1512 VPWR \$3232 \$3200 \$3174 VPWR VGND \$2680 \$3116 VGND
+ sky130_fd_sc_hd__or4_1
X$1513 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1514 VPWR \$3214 VPWR VGND \$2659 VGND sky130_fd_sc_hd__buf_4
X$1515 VPWR \$3200 \$3233 \$2874 VPWR VGND \$2639 \$2837 VGND
+ sky130_fd_sc_hd__or4_1
X$1516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1519 VPWR \$3176 VGND \$3141 VPWR \$1979 VGND sky130_fd_sc_hd__nor2_1
X$1520 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1521 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1526 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1527 VPWR \$2342 \$3305 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1528 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1529 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1530 VPWR \$2780 \$3270 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1531 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1532 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1533 VGND \$856 \$3158 \$2556 \$3202 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$1534 VGND \$856 \$3159 \$2556 \$3215 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$1535 VPWR \$3132 \$3159 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1536 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1538 VPWR \$3031 VGND VPWR \$3216 \$2229 \$3217 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$1539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1540 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1542 VPWR \$1004 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1543 VPWR \$3234 VGND VPWR \$3216 \$2927 \$1004 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$1544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1545 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1546 VGND \$3040 \$3219 \$3017 \$2809 \$3218 \$3131 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1548 VPWR \$3085 VGND VPWR \$3217 \$3143 \$3037 \$2497 VGND
+ sky130_fd_sc_hd__o22a_1
X$1549 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1550 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1551 VGND \$3146 \$3220 \$2403 \$2325 \$3204 \$3262 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1554 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1555 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1556 VGND \$3185 \$3221 \$2971 \$3181 \$3121 \$2880 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1559 VPWR \$3235 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1561 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1562 VPWR \$747 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1565 VGND \$3207 \$2881 \$3236 \$2369 \$2357 \$3004 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1566 VPWR VGND VPWR \$2567 \$3237 \$3398 \$3208 \$3207 VGND
+ sky130_fd_sc_hd__and4_1
X$1567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1568 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1569 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1570 VGND \$3238 \$3108 \$2449 \$2047 \$2048 \$3222 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1571 VGND \$3239 \$1927 \$2005 \$3223 \$3187 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$1572 VPWR \$3240 VGND VPWR \$2360 \$1956 \$3005 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$1573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1574 VGND \$3224 \$3189 \$3225 \$1169 VPWR \$1975 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$1575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1576 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1578 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1579 VGND \$3241 \$3226 \$620 \$1953 \$1987 \$3111 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1581 VGND \$3210 \$3191 \$3242 \$1839 \$2785 \$3038 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1582 VGND \$3192 \$3112 \$2005 \$3227 \$3241 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$1583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1584 VGND \$3211 \$3228 \$2307 \$2180 \$927 \$3194 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1585 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1586 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1587 VGND \$1152 \$3150 \$2450 \$3229 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1589 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1590 VPWR \$3263 \$3138 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1591 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1592 VPWR VGND \$2672 VPWR \$3195 VGND sky130_fd_sc_hd__clkbuf_4
X$1593 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1594 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1595 VPWR VGND \$2694 \$1171 \$3244 \$3212 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1596 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1597 VGND \$2989 \$3244 \$2450 \$3212 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$1598 VGND \$2989 \$3170 \$2232 \$3196 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1599 VPWR VGND \$3169 \$542 \$3213 \$3197 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1601 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1602 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1605 VGND spimemio_flash_clk \$401 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1609 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1611 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1612 VPWR \$5425 VPWR VGND \$5404 \$2472 \$5326 VGND sky130_fd_sc_hd__or3_1
X$1613 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1615 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1616 VGND \$5422 \$4250 \$4892 VPWR VPWR VGND sky130_fd_sc_hd__nand2_4
X$1617 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1618 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1619 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1622 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1623 VPWR \$5304 VGND \$2472 VPWR \$5415 VGND sky130_fd_sc_hd__nor2_1
X$1624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1625 VGND \$5423 \$4617 \$4250 \$4757 \$2741 VPWR VPWR VGND
+ sky130_fd_sc_hd__o31ai_4
X$1626 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1629 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1630 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1631 VPWR VPWR \$5149 VGND \$1315 \$5431 \$5329 VGND sky130_fd_sc_hd__o21ai_1
X$1632 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1633 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1634 VPWR \$5407 VGND \$5184 VPWR \$5532 VGND sky130_fd_sc_hd__nor2_1
X$1635 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1637 VPWR VPWR \$5270 VGND \$1315 \$5426 \$5203 VGND sky130_fd_sc_hd__o21ai_1
X$1638 VPWR VPWR \$5532 VGND \$1315 \$5416 \$5224 VGND sky130_fd_sc_hd__o21ai_1
X$1639 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1641 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1642 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1647 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1649 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1651 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1652 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1653 VPWR VGND \$5252 \$1171 \$5365 \$5409 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1654 VPWR VGND \$5252 \$3694 \$5417 \$5433 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1657 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1660 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1661 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1663 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1664 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1665 VPWR VGND \$5252 \$184 \$5392 \$5410 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1667 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1668 VPWR \$4625 \$5424 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1669 VGND \$4761 \$5424 \$5272 \$5418 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1670 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1671 VPWR VGND \$5332 \$184 \$5419 \$5427 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1673 VPWR VGND VPWR \$3677 \$5419 VGND sky130_fd_sc_hd__inv_2
X$1674 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1675 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1677 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1678 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1681 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1682 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1684 VPWR \$3172 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1685 VGND \$5412 \$3172 \$5385 \$3438 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1686 VGND \$4764 \$5413 \$5298 \$5411 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$1687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1688 VPWR VGND \$5335 \$4774 \$5420 \$5428 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1689 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1692 VGND \$5429 \$4774 \$5420 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$1693 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1694 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1695 VPWR \$5393 VGND VPWR mgmt_gpio_in[17] VGND sky130_fd_sc_hd__clkbuf_1
X$1696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1699 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1700 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1701 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1702 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1703 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1704 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1705 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1706 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1710 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1711 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1714 VPWR \$5434 \$4008 VGND \$5425 \$4807 VPWR VGND sky130_fd_sc_hd__nand3b_1
X$1715 VPWR \$5376 VGND \$5434 \$5440 VPWR VGND sky130_fd_sc_hd__or2_1
X$1716 VPWR VPWR \$5449 VGND \$5326 \$5328 \$5425 VGND sky130_fd_sc_hd__o21ai_1
X$1717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1718 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1719 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1722 VPWR \$5430 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$1723 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1724 VPWR \$5442 VGND VPWR \$5430 VGND sky130_fd_sc_hd__clkbuf_1
X$1725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1726 VPWR \$5435 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$1727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1728 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1729 VPWR \$5443 VGND VPWR \$5435 VGND sky130_fd_sc_hd__clkbuf_1
X$1730 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1731 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1733 VPWR VGND VPWR \$5149 \$5432 VGND sky130_fd_sc_hd__inv_2
X$1734 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1735 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1737 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1740 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1742 VGND \$5436 \$1949 VPWR VPWR VGND sky130_fd_sc_hd__inv_12
X$1743 VPWR \$5097 \$5081 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1745 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1747 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1748 VPWR VGND \$5462 \$2600 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$1749 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1751 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1752 VPWR VGND \$5229 \$411 \$5437 \$5444 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1753 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1754 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1755 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1757 VPWR VGND VPWR \$4278 \$5437 VGND sky130_fd_sc_hd__inv_2
X$1758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1759 VGND \$4761 \$5417 \$4994 \$5433 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1760 VPWR \$2960 \$5417 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$1761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1763 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1768 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1769 VPWR VGND \$5332 \$411 \$5424 \$5418 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1771 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1773 VGND \$4761 \$5419 \$5272 \$5427 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1777 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1778 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1781 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1784 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1785 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1786 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1787 VGND \$4764 \$5420 \$5298 \$5428 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1788 VGND \$4764 \$5454 \$5298 \$5438 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1789 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1790 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1791 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1792 VPWR \$1892 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1793 VPWR \$5446 VGND VPWR \$1892 VGND sky130_fd_sc_hd__clkbuf_1
X$1794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1795 VGND qspi_enabled \$3636 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$1796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1797 VPWR \$3591 VGND VPWR \$3592 \$3531 \$1523 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$1798 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1799 VGND \$3593 \$1897 \$2424 \$3614 \$3322 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$1800 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1801 VGND \$3612 \$3570 \$3409 \$3613 VPWR VPWR \$3067 VGND
+ sky130_fd_sc_hd__or4b_1
X$1802 VPWR \$3613 VPWR VGND \$3483 \$3358 \$3615 VGND sky130_fd_sc_hd__or3b_1
X$1803 VPWR \$2363 \$3570 VGND \$3616 VPWR \$3637 \$1978 VGND
+ sky130_fd_sc_hd__or4_2
X$1804 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1805 VPWR \$3267 VGND \$3617 \$3650 VPWR VGND sky130_fd_sc_hd__or2_1
X$1806 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1808 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1809 VPWR \$3595 VPWR VGND \$3501 \$2640 \$2471 VGND sky130_fd_sc_hd__or3_2
X$1810 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1811 VPWR VGND \$3595 \$2931 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$1812 VPWR \$3596 VGND VPWR \$3452 \$2257 VGND sky130_fd_sc_hd__or2_4
X$1813 VPWR \$3157 \$3618 \$3639 VPWR VGND \$2197 \$3594 VGND
+ sky130_fd_sc_hd__or4_1
X$1814 VPWR \$3442 VGND \$3560 \$3548 VPWR VGND sky130_fd_sc_hd__or2_1
X$1815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1817 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1818 VPWR \$3598 VGND VPWR \$3618 VGND sky130_fd_sc_hd__clkbuf_1
X$1819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1820 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1821 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1824 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1825 VPWR \$2982 \$3668 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1828 VGND \$2777 \$3574 \$3413 \$3619 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1829 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1832 VGND \$856 \$3641 \$3413 \$3640 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1833 VPWR \$3620 VGND \$1059 \$1571 VPWR VGND sky130_fd_sc_hd__or2_1
X$1834 VGND \$3620 \$2474 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$1835 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1836 VPWR \$1570 VGND VPWR \$3204 \$1059 VGND sky130_fd_sc_hd__or2_4
X$1837 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1838 VPWR \$1571 VGND VPWR \$3621 \$1434 VGND sky130_fd_sc_hd__or2_4
X$1839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1843 VPWR \$3576 VGND VPWR \$2464 \$1867 \$3643 \$3562 VGND
+ sky130_fd_sc_hd__o22a_1
X$1844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1845 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1846 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1847 VPWR VGND VPWR \$3578 \$3599 \$3600 \$3622 \$3555 VGND
+ sky130_fd_sc_hd__and4_1
X$1848 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1849 VPWR \$3534 VGND VPWR \$2957 \$3621 \$3623 \$1839 VGND
+ sky130_fd_sc_hd__o22a_1
X$1850 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1852 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1853 VPWR \$3463 VGND VPWR \$3642 \$3621 \$3644 \$1839 VGND
+ sky130_fd_sc_hd__o22a_1
X$1854 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1855 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1858 VPWR \$3602 VGND VPWR \$3645 \$1966 \$2599 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$1859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1860 VPWR \$3582 VGND VPWR \$3624 \$1966 \$3265 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$1861 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1863 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1865 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1866 VPWR \$2431 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1867 VGND \$3626 \$1619 \$3625 \$2649 \$3606 VPWR VPWR VGND
+ sky130_fd_sc_hd__nand4b_4
X$1868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1869 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1870 VPWR \$3625 VPWR VGND \$3607 \$3627 VGND sky130_fd_sc_hd__nand2_1
X$1871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1872 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1873 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1875 VGND \$3646 \$3275 \$2848 \$2047 \$2048 \$3628 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1876 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1877 VPWR \$3647 VGND VPWR \$3294 \$2325 \$3629 \$2918 VGND
+ sky130_fd_sc_hd__o22a_1
X$1878 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1879 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1880 VPWR \$269 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1882 VPWR \$269 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1883 VPWR VGND \$3630 \$1594 \$3546 \$3610 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1884 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1885 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1887 VGND \$2989 \$3589 \$3425 \$3632 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1888 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1889 VGND \$3633 \$3425 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$1890 VPWR VGND VPWR \$3623 \$3529 VGND sky130_fd_sc_hd__inv_2
X$1891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1892 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1893 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1894 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1895 VPWR VGND VPWR \$3644 \$3634 VGND sky130_fd_sc_hd__inv_2
X$1896 VPWR VGND \$3169 \$386 \$3634 \$3635 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1897 VGND \$2989 \$3634 \$3590 \$3635 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$1898 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1901 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1902 VPWR VGND VPWR \$3531 \$3547 VGND sky130_fd_sc_hd__inv_2
X$1903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1904 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1905 VGND \$3322 \$3679 \$3358 \$3661 VPWR VPWR \$3139 VGND
+ sky130_fd_sc_hd__or4b_1
X$1906 VPWR \$3648 \$3649 VGND \$3483 VPWR \$2222 \$3679 VGND
+ sky130_fd_sc_hd__or4_2
X$1907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1908 VPWR \$3650 VPWR VGND \$3614 \$3662 VGND sky130_fd_sc_hd__nand2_1
X$1909 VPWR \$3662 VGND \$3124 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$1910 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1911 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1912 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1913 VGND \$3681 \$3452 \$3471 \$3485 \$3650 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$1914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1916 VPWR VGND VPWR \$3596 \$2700 VGND sky130_fd_sc_hd__inv_2
X$1917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1918 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1919 VPWR \$2197 \$3665 \$3571 VPWR VGND \$3664 \$3663 VGND
+ sky130_fd_sc_hd__or4_1
X$1920 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1923 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1924 VPWR \$3652 VGND \$3572 \$3505 VPWR VGND sky130_fd_sc_hd__or2_1
X$1925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1926 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1927 VPWR \$3682 VGND VPWR \$3665 VGND sky130_fd_sc_hd__clkbuf_1
X$1928 VGND \$1888 \$3666 \$3682 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$1929 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1930 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1931 VPWR VGND \$3667 \$281 \$3668 \$3683 \$3669 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1933 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1934 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1936 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1937 VPWR \$2341 \$3684 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$1938 VPWR VGND \$3670 \$294 \$2877 \$3685 \$3653 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1939 VPWR VGND \$3670 \$281 \$3574 \$3619 \$3653 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1940 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1941 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1942 VPWR VGND \$3435 \$183 \$3641 \$3640 \$3458 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1943 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1944 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1945 VPWR VPWR VGND \$3654 \$3458 VGND sky130_fd_sc_hd__clkbuf_2
X$1946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1947 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1948 VPWR \$3654 VGND \$3143 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$1949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1950 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1953 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1954 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1955 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1960 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1961 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1962 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1963 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1964 VGND \$3671 \$3264 \$2464 \$2047 \$2048 \$3768 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1965 VPWR \$3329 VGND VPWR \$3722 \$2927 \$3444 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$1966 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1968 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1969 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1970 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$1972 VGND \$3421 \$3672 \$553 \$1562 \$2667 \$3673 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1973 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1974 VPWR \$3655 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$1975 VGND \$3605 \$3655 \$3674 \$1219 \$1125 \$3675 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1976 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1977 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1978 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$1979 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1981 VPWR \$3686 VGND VPWR \$1480 \$1776 \$3674 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$1982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$1983 VGND \$3656 \$3676 \$2548 \$1867 \$2667 \$3677 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1984 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1985 VGND \$3687 \$3266 \$2548 \$2047 \$2048 \$3970 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1986 VPWR \$3657 VGND VPWR \$3678 \$1966 \$3465 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$1987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1988 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1989 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$1990 VGND \$3658 \$3647 \$4244 \$2986 \$1867 \$2848 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$1991 VPWR VGND VPWR \$3626 \$3784 \$3659 \$3383 \$3658 VGND
+ sky130_fd_sc_hd__and4_1
X$1992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$1993 VPWR VGND VPWR \$3630 \$3631 VGND sky130_fd_sc_hd__inv_2
X$1994 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1995 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$1996 VPWR VGND \$3630 \$542 \$3589 \$3632 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$1997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$1998 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$1999 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2000 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2001 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2002 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2003 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2005 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2006 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2008 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2009 VGND \$3914 \$3277 \$3953 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$2010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2011 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2012 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2013 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2014 VGND \$2408 \$3593 \$3931 \$3975 \$2537 \$2001 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_2
X$2015 VPWR \$3612 VGND \$3954 \$1897 VPWR VGND sky130_fd_sc_hd__or2_1
X$2016 VPWR VPWR \$3954 VGND \$2815 \$3955 \$3615 VGND sky130_fd_sc_hd__o21ai_1
X$2017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2018 VPWR \$3917 VGND \$3955 \$3956 VPWR VGND sky130_fd_sc_hd__or2_1
X$2019 VGND \$3906 \$3452 \$3471 \$3472 \$3956 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$2020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2021 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2023 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2025 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2026 VPWR \$3976 VGND \$3560 \$3456 VPWR VGND sky130_fd_sc_hd__or2_1
X$2027 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2028 VPWR \$3977 VPWR VGND \$3957 \$3881 VGND sky130_fd_sc_hd__nand2_1
X$2029 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2030 VPWR \$3957 \$3958 VPWR \$2949 VGND \$2741 VGND sky130_fd_sc_hd__o21ba_1
X$2031 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2032 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2034 VGND \$2777 \$3893 \$3413 \$3933 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2037 VPWR VGND VPWR \$3670 \$3653 VGND sky130_fd_sc_hd__inv_2
X$2038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2039 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2040 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2042 VPWR \$3959 VGND \$2366 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$2043 VPWR VPWR VGND \$3959 \$3653 VGND sky130_fd_sc_hd__clkbuf_2
X$2044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2051 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2052 VPWR \$3960 VGND VPWR \$3391 \$2927 \$1076 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$2053 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2054 VGND \$3512 \$3960 \$3961 \$2830 \$2651 \$3910 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2056 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2057 VGND \$3394 \$3962 \$3514 \$2116 \$1536 \$3963 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2058 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2059 VGND \$2160 \$4082 \$2670 \$2646 \$1837 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$2060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2061 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2062 VPWR \$3978 VGND VPWR \$3527 \$2751 \$3961 \$3204 VGND
+ sky130_fd_sc_hd__o22a_1
X$2063 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2064 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2065 VGND \$3795 \$3964 \$1671 \$2809 \$3218 \$3979 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2066 VPWR \$3964 VGND VPWR \$3623 \$2254 \$3581 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$2067 VPWR \$3980 VGND VPWR \$803 \$2724 \$3536 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$2068 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2069 VPWR \$3981 VGND VPWR \$1030 \$2724 \$3965 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$2070 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2071 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2072 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2073 VGND \$3982 \$3981 \$2600 \$2369 \$2357 \$3886 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2076 VGND \$3983 \$3966 \$3967 \$2750 \$2541 \$3292 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2077 VPWR \$3966 VGND VPWR \$3866 \$2559 \$1616 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$2078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2079 VGND \$3984 \$3968 \$3538 \$2116 \$1536 \$1628 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2081 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2082 VPWR \$3985 VGND VPWR \$3885 \$2724 \$2531 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$2083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2085 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2086 VPWR \$3986 VGND VPWR \$925 \$2724 \$3188 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$2087 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2088 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2089 VPWR \$3676 \$3969 VPWR \$3970 VGND \$2581 \$3924 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$2090 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2091 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2092 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2093 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2094 VGND \$3987 \$3971 \$3168 \$2116 \$1536 \$1306 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2096 VGND \$3798 \$3930 \$3899 \$3121 \$2986 \$4145 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2098 VPWR VGND \$3630 \$184 \$3972 \$3988 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2099 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2100 VPWR VGND VPWR \$3292 \$3949 VGND sky130_fd_sc_hd__inv_2
X$2101 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2102 VGND \$2989 \$3949 \$3425 \$3989 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$2103 VGND \$2989 \$3950 \$3590 \$3951 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$2104 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2105 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2106 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2107 VPWR VGND \$3872 \$411 \$3973 \$3990 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2108 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2109 VGND \$2989 \$4005 \$3590 \$3991 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2113 VPWR VGND wb_dat_o[1] VPWR \$3279 VGND sky130_fd_sc_hd__buf_2
X$2114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2115 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2116 VPWR \$3853 \$3699 VPWR \$2336 VGND \$3993 \$3915 VGND
+ sky130_fd_sc_hd__o211ai_1
X$2117 VGND \$3915 \$2336 \$1897 \$3470 \$3833 \$3994 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$2118 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2119 VPWR \$3614 VGND \$3057 \$3994 VPWR VGND sky130_fd_sc_hd__or2_1
X$2120 VPWR \$3615 VGND \$3470 \$3994 VPWR VGND sky130_fd_sc_hd__or2_1
X$2121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2122 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2123 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2126 VGND \$3058 \$3995 \$3124 \$2944 \$2944 \$4049 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2127 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2128 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2129 VPWR \$4007 VGND \$2015 \$4006 VPWR VGND sky130_fd_sc_hd__or2_1
X$2130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2131 VPWR \$3859 VPWR VGND \$3709 \$1998 VGND sky130_fd_sc_hd__or2_2
X$2132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2133 VPWR \$4008 VPWR VGND \$3700 \$3976 VGND sky130_fd_sc_hd__or2_2
X$2134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2135 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2136 VPWR \$3860 VGND \$3710 VPWR \$2815 VGND sky130_fd_sc_hd__nor2_1
X$2137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2138 VPWR \$4009 VGND \$3860 VPWR \$3977 VGND sky130_fd_sc_hd__nor2_1
X$2139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2140 VPWR \$4010 VGND \$2944 VPWR \$2949 VGND sky130_fd_sc_hd__nor2_1
X$2141 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2144 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2145 VPWR VGND \$3667 \$183 \$4012 \$4011 \$3669 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2146 VPWR VGND VPWR \$3667 \$3669 VGND sky130_fd_sc_hd__inv_2
X$2147 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2148 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2150 VPWR \$4013 VGND \$3042 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$2151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2152 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2153 VPWR VGND \$3670 \$183 \$3997 \$3992 \$3653 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2156 VPWR \$3348 \$3996 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2157 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2158 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2159 VPWR VGND VPWR \$2122 \$3997 VGND sky130_fd_sc_hd__inv_2
X$2160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2161 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2163 VPWR VGND VPWR \$2072 \$3998 VGND sky130_fd_sc_hd__inv_2
X$2164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2166 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2168 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2169 VPWR \$3962 VGND \$2007 \$3961 VPWR VGND sky130_fd_sc_hd__or2_1
X$2170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2171 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2172 VGND \$2028 \$3999 \$2670 \$2646 \$3963 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$2173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2174 VGND \$3460 \$3978 \$3575 \$3556 \$3765 \$3943 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2175 VPWR \$3940 VGND VPWR \$3842 \$2927 \$3312 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$2176 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2177 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2178 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2184 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2185 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2186 VPWR VGND VPWR \$3448 \$3942 \$4015 \$3983 \$3982 VGND
+ sky130_fd_sc_hd__and4_1
X$2187 VPWR \$3968 VGND \$2007 \$4039 VPWR VGND sky130_fd_sc_hd__or2_1
X$2188 VPWR VGND VPWR \$4001 \$3941 \$3984 \$3604 \$4016 VGND
+ sky130_fd_sc_hd__and4_1
X$2189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2190 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2192 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2195 VGND \$4018 \$4002 \$3478 \$2750 \$2541 \$3970 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2197 VPWR \$3971 VGND \$2007 \$4017 VPWR VGND sky130_fd_sc_hd__or2_1
X$2198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2199 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2200 VPWR VGND VPWR \$4019 \$3928 \$3987 \$3608 \$4003 VGND
+ sky130_fd_sc_hd__and4_1
X$2201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2202 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2204 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2205 VPWR VGND VPWR \$3970 \$3972 VGND sky130_fd_sc_hd__inv_2
X$2206 VGND \$2989 \$3972 \$4164 \$3988 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2207 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2208 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2209 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2210 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2212 VPWR \$3402 \$4004 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2213 VGND \$2989 \$4004 \$3590 \$4020 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2214 VGND \$2989 \$3973 \$3590 \$3990 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2215 VPWR VGND \$3872 \$386 \$4005 \$3991 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2216 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2217 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2220 VGND \$5280 \$5002 \$5777 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$2221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2222 VPWR \$5755 VGND VPWR \$5302 \$5439 \$5448 \$1975 VGND
+ sky130_fd_sc_hd__o22a_1
X$2223 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2224 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2225 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2226 VPWR VGND \$4853 \$4880 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2227 VPWR VGND VPWR \$4863 \$4891 VGND sky130_fd_sc_hd__inv_2
X$2228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2229 VPWR \$5801 VPWR VGND \$5824 \$5872 \$5778 VGND sky130_fd_sc_hd__or3_1
X$2230 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2231 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2233 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2234 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2236 VPWR \$5779 VGND \$5679 \$5699 VPWR VGND sky130_fd_sc_hd__or2_1
X$2237 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2238 VGND \$5779 \$5770 \$5790 \$5685 VPWR VPWR \$5802 VGND
+ sky130_fd_sc_hd__or4b_1
X$2239 VGND \$5746 \$5648 \$5774 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2241 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2243 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2244 VGND \$5764 \$5791 \$5775 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2245 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2246 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2247 VGND \$5692 \$5792 \$5780 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2249 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2250 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2252 VPWR \$5423 \$5805 VPWR \$5756 VGND VGND sky130_fd_sc_hd__and2_1
X$2253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2254 VGND \$5495 \$5079 \$5803 \$5781 \$5782 \$5765 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2255 VPWR \$5423 \$5781 VPWR \$5783 VGND VGND sky130_fd_sc_hd__and2_1
X$2256 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2257 VGND \$5495 \$5079 \$5749 \$5784 \$5785 \$5786 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2260 VPWR \$5423 \$5806 VPWR \$5787 VGND VGND sky130_fd_sc_hd__and2_1
X$2261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2262 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2263 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2265 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2266 VPWR VGND \$5559 \$3711 \$5750 \$5807 \$5553 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2268 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2270 VPWR VGND \$5388 \$1171 \$5751 \$5808 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2272 VPWR VGND \$5388 \$3694 \$5776 \$5809 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2273 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2274 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2277 VGND \$2777 \$5793 \$5408 \$5771 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$2278 VPWR VGND \$5525 \$3694 \$5793 \$5771 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2279 VPWR VGND VPWR \$5788 \$1615 VGND sky130_fd_sc_hd__inv_4
X$2280 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2281 VPWR VGND \$5525 \$3711 \$5752 \$5757 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2282 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2283 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2285 VGND \$5528 \$2854 mgmt_gpio_out[20] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2286 VPWR \$5810 VGND VPWR \$2111 VGND sky130_fd_sc_hd__clkbuf_1
X$2287 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2289 VPWR \$5811 VGND VPWR \$2960 VGND sky130_fd_sc_hd__clkbuf_1
X$2290 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2291 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2294 VGND \$5413 \$2960 mgmt_gpio_out[23] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2295 VPWR \$5796 VGND VPWR \$1320 VGND sky130_fd_sc_hd__clkbuf_1
X$2296 VGND \$4761 \$5730 \$5272 \$5738 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2297 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2298 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2299 VPWR \$5797 VGND VPWR \$5789 VGND sky130_fd_sc_hd__clkbuf_1
X$2300 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2301 VPWR \$5772 VGND VPWR \$1373 VGND sky130_fd_sc_hd__clkbuf_1
X$2302 VGND \$4761 \$5758 \$5334 \$5767 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2303 VGND \$4761 \$5759 \$5334 \$5742 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2304 VPWR \$5798 VGND VPWR \$1949 VGND sky130_fd_sc_hd__clkbuf_1
X$2305 VPWR \$5773 VGND VPWR \$1221 VGND sky130_fd_sc_hd__clkbuf_1
X$2306 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2308 VGND \$4764 \$5760 \$5334 \$5768 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2309 VGND \$4764 \$5731 \$5298 \$5739 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$2310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2311 VPWR \$5812 VGND VPWR \$5904 VGND sky130_fd_sc_hd__clkbuf_1
X$2312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2313 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2316 VGND \$5732 \$1023 mgmt_gpio_out[19] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2319 VPWR VPWR VGND spimemio_flash_io2_oeb \$5870 VGND
+ sky130_fd_sc_hd__clkbuf_2
X$2320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2321 VGND \$5777 \$5280 \$5439 \$2221 \$5448 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$2322 VPWR VGND \$5823 VPWR spimemio_flash_io3_do VGND
+ sky130_fd_sc_hd__clkbuf_4
X$2323 VPWR \$5882 VGND VPWR \$5616 VGND sky130_fd_sc_hd__clkbuf_1
X$2324 VPWR \$4833 \$4864 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$2325 VGND \$5873 \$4833 \$5872 \$5824 \$4863 VPWR VPWR VGND
+ sky130_fd_sc_hd__nand4bb_1
X$2326 VPWR \$5824 VGND VPWR wb_adr_i[9] VGND sky130_fd_sc_hd__clkbuf_1
X$2327 VPWR \$5841 \$5778 \$5813 VPWR VGND \$5834 \$5840 VGND
+ sky130_fd_sc_hd__or4_1
X$2328 VPWR \$4880 \$5715 \$5814 VPWR VGND \$5897 \$5873 VGND
+ sky130_fd_sc_hd__or4_1
X$2329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2330 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2331 VPWR \$5814 VPWR VGND \$5842 \$5815 VGND sky130_fd_sc_hd__nand2_1
X$2332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2333 VPWR \$5842 \$5883 \$5815 VPWR VGND \$5825 \$5835 VGND
+ sky130_fd_sc_hd__or4_1
X$2334 VPWR \$5843 VPWR \$5825 \$5745 \$5835 \$5875 VGND VGND
+ sky130_fd_sc_hd__nand4_1
X$2335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2336 VPWR \$5659 VGND \$5684 \$5458 VPWR \$5779 VGND sky130_fd_sc_hd__o21ai_2
X$2337 VGND \$5471 \$5659 \$5684 \$5779 \$5685 \$5836 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$2338 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2339 VPWR \$5836 VPWR VGND \$5845 \$5844 VGND sky130_fd_sc_hd__nand2_1
X$2340 VGND \$5876 \$5884 \$5846 \$5875 VPWR VPWR \$5843 VGND
+ sky130_fd_sc_hd__or4b_1
X$2341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2342 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2344 VGND \$5802 \$5847 \$5848 \$5849 VPWR VPWR \$5816 VGND
+ sky130_fd_sc_hd__or4bb_1
X$2345 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2346 VPWR \$5877 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2347 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2348 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2349 VPWR \$5877 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2350 VGND \$5790 \$5837 \$5877 \$5850 VPWR VPWR \$5817 VGND
+ sky130_fd_sc_hd__or4bb_1
X$2351 VGND \$5774 \$5885 \$5804 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2353 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2354 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2355 VGND \$5691 \$5886 \$5851 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2356 VGND \$5729 \$5826 \$5749 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2357 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2358 VGND \$5717 \$5934 \$5818 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2359 VGND \$5495 \$5079 \$5818 \$5805 \$5852 \$5853 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2360 VGND \$5495 \$5079 \$5804 \$5854 \$5935 \$5855 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2361 VGND \$5495 \$5079 \$5851 \$5819 \$5936 \$5856 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2362 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2363 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2364 VGND \$5495 \$5079 \$5775 \$5857 \$5878 \$5858 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2365 VGND \$5495 \$5079 \$5780 \$5806 \$5827 \$5859 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$2366 VPWR \$5423 \$5819 VPWR \$5860 VGND VGND sky130_fd_sc_hd__and2_1
X$2367 VPWR \$5423 \$5857 VPWR \$5861 VGND VGND sky130_fd_sc_hd__and2_1
X$2368 VPWR \$5423 \$5784 VPWR \$5862 VGND VGND sky130_fd_sc_hd__and2_1
X$2369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2370 VGND \$2777 \$5750 \$5165 \$5807 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$2371 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2372 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2373 VGND \$2777 \$5751 \$5408 \$5808 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$2374 VGND \$2777 \$5776 \$5408 \$5809 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$2375 VPWR \$4584 \$5776 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$2376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2377 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2378 VGND \$2111 \$5793 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$2379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2380 VPWR \$3122 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2381 VGND \$5887 \$3122 \$5870 \$3636 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$2382 VPWR \$4230 \$5863 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2384 VPWR \$5879 VGND VPWR \$2854 VGND sky130_fd_sc_hd__clkbuf_1
X$2385 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2386 VPWR \$5888 VGND VPWR \$5879 VGND sky130_fd_sc_hd__clkbuf_1
X$2387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2388 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2389 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2391 VPWR \$5889 VGND VPWR \$5864 VGND sky130_fd_sc_hd__clkbuf_1
X$2392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2393 VPWR \$5864 VGND VPWR \$1821 VGND sky130_fd_sc_hd__clkbuf_1
X$2394 VGND \$5652 \$2111 mgmt_gpio_out[22] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2395 VGND \$5731 \$1821 mgmt_gpio_out[21] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2396 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2397 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2398 VGND \$5730 \$3037 mgmt_gpio_out[24] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2399 VPWR VGND \$5865 \$3136 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2400 VPWR \$5890 VGND VPWR \$1925 VGND sky130_fd_sc_hd__clkbuf_1
X$2401 VPWR \$5789 VGND VPWR \$500 VGND sky130_fd_sc_hd__clkbuf_1
X$2402 VGND \$5758 \$500 mgmt_gpio_out[27] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2403 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2404 VPWR \$5831 VGND VPWR \$5772 VGND sky130_fd_sc_hd__clkbuf_1
X$2405 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2406 VGND \$5759 \$1855 mgmt_gpio_out[29] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2407 VPWR VGND VPWR \$5008 \$5866 VGND sky130_fd_sc_hd__inv_2
X$2408 VGND \$5832 \$5733 \$5658 \$3636 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2409 VPWR \$5891 VGND VPWR \$5773 VGND sky130_fd_sc_hd__clkbuf_1
X$2410 VPWR \$5880 VGND VPWR \$4584 VGND sky130_fd_sc_hd__clkbuf_1
X$2411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2412 VPWR \$5892 VGND VPWR \$5880 VGND sky130_fd_sc_hd__clkbuf_1
X$2413 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2414 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2416 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2417 VPWR \$5893 VGND VPWR \$5769 VGND sky130_fd_sc_hd__clkbuf_1
X$2418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2419 VGND \$5760 \$3092 mgmt_gpio_out[34] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2420 VPWR VGND \$5867 \$3137 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2422 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2423 VPWR \$5753 VGND VPWR mgmt_gpio_in[19] VGND sky130_fd_sc_hd__clkbuf_1
X$2424 VPWR \$5894 VGND VPWR \$5868 VGND sky130_fd_sc_hd__clkbuf_1
X$2425 VPWR \$5868 VGND VPWR \$1023 VGND sky130_fd_sc_hd__clkbuf_1
X$2426 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2427 VPWR VGND mgmt_gpio_out[37] VPWR \$5929 VGND sky130_fd_sc_hd__buf_2
X$2428 VPWR VGND mgmt_gpio_out[36] VPWR \$5832 VGND sky130_fd_sc_hd__buf_2
X$2429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2432 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2433 VPWR \$311 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2434 VPWR \$311 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2435 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2436 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2438 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2439 VPWR \$5633 VPWR \$5647 VGND \$4880 \$5147 VGND sky130_fd_sc_hd__o21a_1
X$2440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2444 VPWR \$5520 VGND VPWR \$5684 \$5682 \$5679 \$5690 VGND
+ sky130_fd_sc_hd__o22a_1
X$2445 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2446 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2448 VGND \$4444 \$5685 \$5684 \$5699 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$2449 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2453 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2455 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2458 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2459 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2462 VPWR \$5613 \$5687 VPWR \$5701 VGND VGND sky130_fd_sc_hd__and2_1
X$2463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2465 VPWR VGND \$5702 \$2524 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2466 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2468 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2469 VPWR VGND \$5559 \$1594 \$5689 \$5710 \$5553 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2470 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2477 VPWR VGND VPWR \$5229 \$5207 VGND sky130_fd_sc_hd__inv_2
X$2478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2481 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2482 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2484 VPWR VGND VPWR \$4053 \$5703 VGND sky130_fd_sc_hd__inv_2
X$2485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2488 VPWR VGND VPWR \$3447 \$5704 VGND sky130_fd_sc_hd__inv_2
X$2489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2491 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2492 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2496 VPWR VGND VPWR \$5705 \$4562 VGND sky130_fd_sc_hd__inv_4
X$2497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2498 VPWR VGND \$5627 \$3711 \$5697 \$5706 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2499 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2500 VGND \$4761 \$5697 \$5272 \$5706 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2502 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2503 VPWR VGND \$5627 \$411 \$5698 \$5694 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2505 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2506 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2511 VGND \$5707 \$184 \$5665 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2513 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2520 VGND spimemio_flash_io1_oeb \$311 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$2521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2523 VPWR \$4733 \$4881 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$2524 VPWR VGND VPWR \$5147 \$4916 VGND sky130_fd_sc_hd__inv_2
X$2525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2526 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2527 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2528 VPWR \$5468 VPWR VGND \$5633 \$4863 \$4833 VGND sky130_fd_sc_hd__or3_2
X$2529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2530 VPWR \$4733 \$5683 \$5274 VPWR VGND \$5745 \$5715 VGND
+ sky130_fd_sc_hd__or4_1
X$2531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2535 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2536 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2537 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2539 VPWR \$5700 VGND VPWR \$5708 VGND sky130_fd_sc_hd__clkbuf_1
X$2540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2542 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2545 VPWR \$5693 VGND VPWR \$5709 VGND sky130_fd_sc_hd__clkbuf_1
X$2546 VGND \$5709 \$5681 \$5717 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2548 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2550 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2552 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2553 VGND \$2777 \$5689 \$5165 \$5710 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2554 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2555 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2556 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2557 VPWR VGND \$5718 \$3035 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2559 VPWR VGND VPWR \$3395 \$5725 VGND sky130_fd_sc_hd__inv_2
X$2560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2561 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2562 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2563 VPWR VGND \$5229 \$3694 \$5720 \$5719 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2566 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2567 VGND \$5720 \$1373 VPWR VPWR VGND sky130_fd_sc_hd__inv_8
X$2568 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2569 VPWR \$1601 \$5711 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$2570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2571 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2572 VGND \$2777 \$5703 \$5367 \$5721 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2573 VPWR VGND VPWR \$4315 \$5712 VGND sky130_fd_sc_hd__inv_2
X$2574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2576 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2577 VGND \$4761 \$5704 \$5367 \$5713 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2578 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2580 VPWR VGND VPWR \$5562 \$5527 VGND sky130_fd_sc_hd__inv_2
X$2581 VPWR VGND \$5562 \$3694 \$5705 \$5714 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2582 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2583 VGND \$4761 \$5705 \$5369 \$5714 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2588 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2592 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2593 VPWR VGND \$5345 \$184 \$5722 \$5723 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2594 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2595 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2596 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2597 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2603 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2604 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2605 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2610 VPWR \$4817 VGND VPWR \$4696 \$4508 \$1619 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$2611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2612 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2613 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2614 VPWR \$3993 VPWR VGND \$3470 \$1979 VGND sky130_fd_sc_hd__or2_2
X$2615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2617 VPWR VPWR \$3993 \$4799 \$4211 \$4602 \$1962 \$3470 VGND VGND
+ sky130_fd_sc_hd__o2111ai_1
X$2618 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2619 VPWR VGND VPWR \$4646 \$4474 VGND sky130_fd_sc_hd__inv_2
X$2620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2621 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2622 VGND \$4786 \$3742 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$2623 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2624 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2626 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2627 VPWR VGND VPWR \$4663 \$4035 VGND sky130_fd_sc_hd__inv_2
X$2628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2630 VPWR \$4370 VPWR VGND \$4772 \$4800 VGND sky130_fd_sc_hd__or2_2
X$2631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2632 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2633 VPWR \$4801 VGND \$4808 \$4736 VPWR VGND sky130_fd_sc_hd__or2_1
X$2634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2635 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2636 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2638 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2639 VPWR \$4788 VPWR VGND \$4758 \$4739 \$4801 VGND sky130_fd_sc_hd__or3_1
X$2640 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2641 VPWR \$4789 VGND \$4788 \$4665 VPWR VGND sky130_fd_sc_hd__or2_1
X$2642 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2643 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2644 VGND \$4774 \$293 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$2645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2646 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2647 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2648 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2649 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2650 VPWR VGND \$4701 \$3711 \$4790 \$4802 \$4677 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2651 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2652 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2654 VPWR VGND \$4803 VPWR \$4791 VGND sky130_fd_sc_hd__clkbuf_4
X$2655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2656 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2660 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2661 VPWR VGND \$4654 \$184 \$4792 \$4804 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2663 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2664 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2665 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2666 VPWR VGND VPWR \$3465 \$4792 VGND sky130_fd_sc_hd__inv_2
X$2667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2671 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2678 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2681 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2682 VGND \$4353 \$4784 \$4765 \$4793 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2683 VPWR VGND VPWR \$4681 \$4682 VGND sky130_fd_sc_hd__inv_2
X$2684 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2685 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2688 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2689 VPWR \$4243 \$4796 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2690 VPWR VGND \$4709 \$411 \$4796 \$4814 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2693 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2694 VPWR VGND \$4805 \$2992 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2696 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2697 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2699 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2701 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2702 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2703 VGND \$4746 mgmt_gpio_in[14] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$2704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2706 VPWR VGND wb_dat_o[17] VPWR \$4816 VGND sky130_fd_sc_hd__buf_2
X$2707 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2708 VGND \$4696 \$4651 \$4817 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$2709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2711 VGND \$3832 \$4615 \$4818 \$4799 \$4806 \$4646 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$2712 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2713 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2714 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2718 VPWR \$4734 VPWR VGND \$2741 \$4035 \$4603 VGND sky130_fd_sc_hd__or3_1
X$2719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2720 VPWR VGND VPWR \$4597 \$1962 VGND sky130_fd_sc_hd__inv_2
X$2721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2722 VPWR \$2336 VPWR VGND \$4807 \$3342 \$4035 VGND sky130_fd_sc_hd__or3_2
X$2723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2724 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2725 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2726 VPWR VPWR \$4673 VGND \$1962 \$4808 \$4834 VGND sky130_fd_sc_hd__o21ai_1
X$2727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2728 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2729 VPWR \$4131 VPWR VGND \$4835 \$4989 VGND sky130_fd_sc_hd__or2_2
X$2730 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2731 VPWR \$4809 VGND \$4787 \$4819 VPWR VGND sky130_fd_sc_hd__or2_1
X$2732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2733 VPWR \$4810 VGND \$4553 \$4809 VPWR VGND sky130_fd_sc_hd__or2_1
X$2734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2735 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2736 VPWR \$4820 VGND \$4572 \$4810 VPWR VGND sky130_fd_sc_hd__or2_1
X$2737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2738 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2740 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2741 VGND \$2777 \$4780 \$4811 \$4812 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2743 VGND \$2777 \$4790 \$4811 \$4802 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$2744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2745 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2749 VPWR VGND VPWR \$3131 \$4836 VGND sky130_fd_sc_hd__inv_2
X$2750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2753 VPWR \$3575 \$4821 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2754 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2755 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2757 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2758 VPWR VGND VPWR \$2784 \$4822 VGND sky130_fd_sc_hd__inv_2
X$2759 VGND \$4761 \$4792 \$4813 \$4804 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2763 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2768 VPWR VGND VPWR \$2547 \$4824 VGND sky130_fd_sc_hd__inv_2
X$2769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2770 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2772 VPWR \$3538 \$4823 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2774 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2775 VGND \$4764 \$4838 \$4850 \$4825 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2779 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2780 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2781 VPWR VPWR VGND \$4783 \$3952 VGND sky130_fd_sc_hd__clkbuf_2
X$2782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2784 VPWR VGND \$4681 \$354 \$4827 \$4826 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2785 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2786 VPWR \$3586 \$4827 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2789 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2790 VGND \$4353 \$4796 \$4427 \$4814 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2792 VPWR VGND \$4709 \$1594 \$4805 \$4815 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2793 VGND \$4353 \$4805 \$4828 \$4815 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2794 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2795 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2796 VGND \$4829 \$4750 \$1171 \$4686 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2798 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2799 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2800 VGND \$4769 \$184 \$4830 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2803 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2805 VPWR \$4832 VGND VPWR \$4831 VGND sky130_fd_sc_hd__clkbuf_1
X$2806 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2807 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2808 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2811 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2812 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2813 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2816 VPWR \$3878 \$3891 \$4456 VPWR VGND \$3906 \$3681 VGND
+ sky130_fd_sc_hd__or4_1
X$2817 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2818 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2819 VPWR \$3892 \$3836 VPWR \$2815 VGND VGND sky130_fd_sc_hd__and2_1
X$2820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2821 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2823 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2824 VPWR \$3907 \$3701 VPWR \$2996 VGND \$3709 VGND sky130_fd_sc_hd__o21ba_1
X$2825 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2828 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2829 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2831 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2833 VPWR VGND VPWR \$3333 \$3893 VGND sky130_fd_sc_hd__inv_2
X$2834 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2835 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2836 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2837 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2842 VPWR VGND \$3894 \$293 \$3895 \$3909 \$3908 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2844 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2845 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2846 VPWR \$2281 \$3895 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$2847 VPWR \$3896 VGND VPWR \$3840 \$2927 \$815 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$2848 VGND \$2721 \$3896 \$3897 \$2830 \$2651 \$3883 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2850 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2851 VPWR \$3911 VGND \$2007 \$3897 VPWR VGND sky130_fd_sc_hd__or2_1
X$2852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2853 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2854 VPWR \$2517 VGND VPWR \$3898 \$2670 \$3934 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$2855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2856 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2857 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2858 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2860 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2861 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2862 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2863 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2868 VPWR \$3750 VGND \$2007 \$3899 VPWR VGND sky130_fd_sc_hd__or2_1
X$2869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2870 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2871 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2872 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2874 VPWR VGND VPWR \$3751 \$3903 \$3902 \$3900 \$3901 VGND
+ sky130_fd_sc_hd__and4_1
X$2875 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2876 VPWR \$3904 VGND \$2007 \$3825 VPWR VGND sky130_fd_sc_hd__or2_1
X$2877 VGND \$3912 \$3904 \$1893 \$2116 \$1536 \$1702 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2878 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2879 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2880 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2881 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2883 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2884 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2886 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2887 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2888 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2889 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2891 VPWR VGND \$3950 \$1616 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2894 VPWR VGND \$3888 \$1671 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$2895 VPWR VGND \$3716 \$1171 \$3888 \$3876 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2896 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2897 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2898 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2901 VGND \$3889 \$2846 mgmt_gpio_out[10] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$2902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2903 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2904 VPWR VGND wb_dat_o[0] VPWR \$3592 VGND sky130_fd_sc_hd__buf_2
X$2905 VPWR \$3953 VGND VPWR \$3914 \$3531 \$2057 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$2906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2908 VGND \$3931 \$3915 \$3612 \$3615 \$3916 \$2001 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$2909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2911 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2912 VGND \$3741 \$3617 \$3918 \$3689 VPWR VPWR \$3917 VGND
+ sky130_fd_sc_hd__or4b_1
X$2913 VGND \$3878 \$3452 \$3471 \$3484 \$3955 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$2914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2916 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2917 VPWR \$3859 \$3919 VPWR \$3907 VGND VGND sky130_fd_sc_hd__and2_1
X$2918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2920 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2921 VPWR VPWR \$3710 VGND \$2931 \$3932 \$3809 VGND sky130_fd_sc_hd__o21bai_1
X$2922 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2925 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2926 VPWR VGND \$3667 \$200 \$3893 \$3933 \$3669 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2929 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2930 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2933 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2934 VGND \$856 \$3884 \$3413 \$3920 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2935 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2936 VPWR VGND \$3894 \$3732 \$3884 \$3920 \$3908 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2937 VGND \$856 \$3895 \$3921 \$3909 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$2938 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2939 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2940 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2941 VPWR \$3922 VGND \$2007 \$3734 VPWR VGND sky130_fd_sc_hd__or2_1
X$2942 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2943 VGND \$3922 \$2685 \$2116 \$1536 \$3934 \$2283 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$2944 VGND \$2860 \$3911 \$2896 \$2116 \$1536 \$3935 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2945 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2946 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2947 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2948 VPWR \$2368 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2949 VGND \$2803 \$2368 \$3936 \$1845 \$2375 \$3937 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2950 VPWR \$3938 VGND VPWR \$1242 \$2724 \$3937 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$2951 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2952 VPWR \$2500 VGND VPWR \$3939 \$2670 \$3935 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$2953 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2954 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2955 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2956 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2957 VGND \$3941 \$3462 \$3923 \$1715 \$1754 \$803 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2959 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2960 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2961 VGND \$3942 \$3940 \$3899 \$2830 \$2651 \$3524 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2962 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2963 VPWR \$3223 VGND VPWR \$3943 \$2670 \$1628 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$2964 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2965 VPWR \$2351 VPWR \$3925 \$4232 \$3924 VGND \$1335 VGND
+ sky130_fd_sc_hd__a22oi_1
X$2966 VGND \$3902 \$3925 \$3885 \$859 \$2789 \$3926 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2967 VGND \$3945 \$3726 \$3926 \$1715 \$1754 \$3885 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2968 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2969 VPWR VGND VPWR \$3947 \$3945 \$3912 \$3516 \$3946 VGND
+ sky130_fd_sc_hd__and4_1
X$2970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2971 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2972 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2973 VGND \$3928 \$3379 \$3927 \$1715 \$1754 \$925 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$2974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$2977 VPWR \$3227 VGND VPWR \$3929 \$2670 \$1306 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$2978 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2979 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2980 VPWR \$826 VPWR \$3930 \$3948 \$3611 VGND \$1335 VGND
+ sky130_fd_sc_hd__a22oi_1
X$2981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2983 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2984 VPWR VGND \$3630 \$1179 \$3949 \$3989 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2987 VPWR VGND \$3716 \$1179 \$3950 \$3951 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$2988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2989 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$2992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$2993 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$2994 VGND \$3952 \$3590 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$2995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$2996 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$2997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$2998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$2999 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3002 VPWR VPWR \$3057 VGND \$2234 \$4033 \$3614 VGND sky130_fd_sc_hd__o21ai_1
X$3003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3004 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3005 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3008 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3010 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3011 VPWR VGND \$3124 VPWR \$4022 VGND sky130_fd_sc_hd__clkbuf_4
X$3012 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3013 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3015 VGND \$4007 \$2234 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$3016 VPWR VGND \$2949 VPWR \$4063 VGND sky130_fd_sc_hd__clkbuf_4
X$3017 VPWR \$2336 \$3560 VGND \$4035 VPWR \$4006 VGND sky130_fd_sc_hd__nor3_1
X$3018 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3019 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3023 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3024 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3025 VGND \$2777 \$4012 \$3413 \$4011 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3026 VPWR VPWR VGND \$4013 \$3669 VGND sky130_fd_sc_hd__clkbuf_2
X$3027 VPWR VGND \$3670 \$200 \$3996 \$4036 \$3653 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3028 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3029 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3030 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3031 VGND \$2777 \$3997 \$3413 \$3992 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3032 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3033 VGND \$4023 \$183 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$3034 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3035 VPWR \$4024 VGND \$3106 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$3036 VPWR VPWR VGND \$4024 \$3908 VGND sky130_fd_sc_hd__clkbuf_2
X$3037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3038 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3039 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3040 VPWR \$4037 VGND VPWR \$3349 \$3106 \$3509 \$3271 VGND
+ sky130_fd_sc_hd__o22a_1
X$3041 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3046 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3047 VPWR \$4038 VGND VPWR \$2122 \$2366 \$3721 \$2751 VGND
+ sky130_fd_sc_hd__o22a_1
X$3048 VGND \$4026 \$4040 \$4025 \$4014 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$3049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3050 VGND \$4026 \$4000 \$3348 \$2366 \$2986 \$4027 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3051 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3052 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3053 VGND \$4014 \$4037 \$3222 \$2581 \$2918 \$4028 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3055 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3056 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3057 VGND \$4041 \$4097 \$4039 \$2830 \$2651 \$3644 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3058 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3062 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3063 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3067 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3068 VPWR \$3887 VGND VPWR \$4029 \$2927 \$3674 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$3069 VGND \$4042 \$3986 \$1099 \$2369 \$2357 \$4030 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3071 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3072 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3073 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3074 VPWR \$4002 VGND VPWR \$4031 \$2559 \$3519 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$3075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3076 VPWR \$4043 VGND VPWR \$3242 \$2254 \$3929 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$3077 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3079 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3080 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3084 VPWR VGND \$3716 \$411 \$4004 \$4020 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3086 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3087 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3088 VPWR \$3541 \$3973 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3090 VPWR \$3943 \$4005 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3092 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3093 VGND mgmt_gpio_in[11] \$1424 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$3094 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3095 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3096 VPWR VGND wb_dat_o[2] VPWR \$3740 VGND sky130_fd_sc_hd__buf_2
X$3097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3099 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3101 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3102 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3103 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3104 VGND \$3691 \$4048 \$4049 \$2931 \$3742 \$2742 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3105 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3106 VPWR \$3029 VGND \$4050 \$4044 VPWR VGND sky130_fd_sc_hd__or2_1
X$3107 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3108 VPWR \$3280 VGND \$4050 \$4077 VPWR VGND sky130_fd_sc_hd__or2_1
X$3109 VPWR \$3214 VGND \$4050 \$4062 VPWR VGND sky130_fd_sc_hd__or2_1
X$3110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3111 VPWR \$3709 VPWR VGND \$2336 \$4035 VGND sky130_fd_sc_hd__or2_2
X$3112 VPWR \$2336 \$3700 VGND \$4035 VPWR \$1979 VGND sky130_fd_sc_hd__nor3_1
X$3113 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3114 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3115 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3118 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3120 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3121 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3123 VGND \$2777 \$3996 \$3413 \$4036 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3126 VGND \$856 \$3998 \$3413 \$4051 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3128 VPWR VGND VPWR \$3894 \$3908 VGND sky130_fd_sc_hd__inv_2
X$3129 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3130 VPWR VGND \$3894 \$3711 \$4046 \$4045 \$3908 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3131 VGND \$856 \$4046 \$3921 \$4045 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3132 VPWR \$2999 \$4064 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3133 VPWR VGND VPWR \$3349 \$4046 VGND sky130_fd_sc_hd__inv_2
X$3134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3135 VGND \$2878 \$4052 \$2783 \$2809 \$3218 \$2597 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3136 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3137 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3138 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3141 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3143 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3144 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3147 VGND \$4047 \$3980 \$3417 \$2369 \$2357 \$4028 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3150 VGND \$4055 \$4054 \$4053 \$2750 \$2541 \$3222 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3151 VGND \$4055 \$4221 \$3252 \$4047 \$4041 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$3152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3154 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3157 VPWR \$4056 VGND VPWR \$3644 \$2254 \$3943 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$3158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3160 VPWR \$4057 VGND VPWR \$4058 \$2927 \$3714 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$3161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3162 VPWR \$3871 VGND VPWR \$4058 \$3019 \$3543 \$2751 VGND
+ sky130_fd_sc_hd__o22a_1
X$3163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3164 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3165 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3166 VPWR \$4059 VGND VPWR \$1856 \$2254 \$3541 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$3167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3170 VGND \$4060 \$4069 \$4017 \$2830 \$2651 \$3242 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3171 VGND \$4018 \$4172 \$3193 \$4042 \$4060 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$3172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3173 VGND \$4003 \$4043 \$3519 \$2809 \$3218 \$4187 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3174 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3175 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3176 VPWR \$3228 VGND VPWR \$4187 \$2921 \$4017 \$3121 VGND
+ sky130_fd_sc_hd__o22a_1
X$3177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3181 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3188 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3194 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3195 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3197 VGND \$4842 \$3470 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_8
X$3198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3200 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3201 VPWR \$4576 VPWR VGND \$4076 \$4833 \$4854 VGND sky130_fd_sc_hd__or3_2
X$3202 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3203 VPWR \$4214 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3204 VPWR \$4214 VPWR VGND \$4044 \$4864 \$4892 VGND sky130_fd_sc_hd__or3_2
X$3205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3207 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3208 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3209 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3210 VPWR VGND VPWR \$4855 \$4734 VGND sky130_fd_sc_hd__inv_2
X$3211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3212 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3213 VPWR \$4834 \$4843 VPWR \$1979 VGND \$4673 VGND sky130_fd_sc_hd__o21ba_1
X$3214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3215 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3216 VPWR \$4835 VGND \$5106 \$4326 VPWR VGND sky130_fd_sc_hd__or2_1
X$3217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3218 VPWR \$4856 VGND \$4835 \$4373 VPWR VGND sky130_fd_sc_hd__or2_1
X$3219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3220 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3222 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3223 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3227 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3228 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3229 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3230 VGND \$2777 \$4836 \$4811 \$4844 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3231 VPWR VGND \$4760 \$3694 \$4836 \$4844 \$4717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3233 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3234 VPWR VGND VPWR \$3537 \$4845 VGND sky130_fd_sc_hd__inv_2
X$3235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3236 VPWR VGND \$4781 \$3711 \$4821 \$4871 \$4782 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3237 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3238 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3239 VGND \$4761 \$4822 \$4813 \$4846 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3240 VPWR VGND \$4654 \$4023 \$4822 \$4846 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3242 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3244 VPWR VGND VPWR \$4237 \$4847 VGND sky130_fd_sc_hd__inv_2
X$3245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3246 VPWR \$3368 \$4848 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3247 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3248 VGND \$4353 \$4857 \$4813 \$4849 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3249 VPWR VGND VPWR \$4274 \$4851 VGND sky130_fd_sc_hd__inv_2
X$3250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3251 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3252 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3253 VPWR VGND \$4681 \$3711 \$4823 \$4837 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3254 VGND \$4764 \$4823 \$4850 \$4837 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3255 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3256 VPWR VGND \$4707 \$411 \$4838 \$4825 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3257 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3258 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3259 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3260 VPWR VGND VPWR \$3926 \$4838 VGND sky130_fd_sc_hd__inv_2
X$3261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3262 VPWR VGND VPWR \$4707 \$4706 VGND sky130_fd_sc_hd__inv_2
X$3263 VPWR VGND \$4707 \$354 \$4839 \$4875 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3265 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3266 VPWR \$3752 \$4839 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3268 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3269 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3270 VGND \$4353 \$4827 \$4427 \$4826 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3273 VPWR VGND \$4709 \$386 \$4840 \$4858 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3274 VPWR VGND VPWR \$4027 \$4840 VGND sky130_fd_sc_hd__inv_2
X$3275 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3276 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3277 VPWR \$4709 \$4710 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3279 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3280 VPWR \$4841 VGND VPWR \$4829 VGND sky130_fd_sc_hd__clkbuf_1
X$3281 VGND \$2989 \$4750 \$4828 \$4841 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$3282 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3283 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3284 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3285 VPWR VGND \$4650 \$184 \$4830 \$4859 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3286 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3287 VGND \$2989 \$3890 \$4828 \$4860 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$3288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3290 VPWR VGND wb_dat_o[18] VPWR \$4862 VGND sky130_fd_sc_hd__buf_2
X$3291 VGND \$4879 \$4601 \$4508 \$4509 \$2221 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$3292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3294 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3295 VGND \$4853 \$2964 \$4863 \$4733 \$4833 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$3296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3298 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3299 VGND \$4733 \$3230 \$4864 \$4853 \$4863 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$3300 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3301 VGND \$4854 \$4864 \$3485 \$4576 VPWR VPWR VGND sky130_fd_sc_hd__nor3_4
X$3302 VPWR VGND \$4035 VPWR \$4902 VGND sky130_fd_sc_hd__clkbuf_4
X$3303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3306 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3307 VPWR \$4865 VGND \$2741 \$4673 VPWR VGND sky130_fd_sc_hd__or2_1
X$3308 VPWR \$4843 VPWR VGND \$4865 \$4903 VGND sky130_fd_sc_hd__nand2_1
X$3309 VPWR VGND VPWR \$4267 \$4865 VGND sky130_fd_sc_hd__inv_2
X$3310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3311 VPWR \$4675 VGND \$4819 \$4866 VPWR VGND sky130_fd_sc_hd__or2_1
X$3312 VPWR \$4487 VGND \$4819 \$4883 VPWR VGND sky130_fd_sc_hd__or2_1
X$3313 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3314 VPWR \$4867 VGND \$4856 \$4882 VPWR VGND sky130_fd_sc_hd__or2_1
X$3315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3316 VPWR \$4884 VPWR VGND \$4739 \$4676 \$4867 VGND sky130_fd_sc_hd__or3_1
X$3317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3318 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3319 VPWR \$4868 VGND \$4885 \$4617 VPWR VGND sky130_fd_sc_hd__or2_1
X$3320 VPWR \$4885 VGND \$4605 VPWR \$4884 VGND sky130_fd_sc_hd__nor2_1
X$3321 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3322 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3323 VPWR \$4869 VGND \$4886 VPWR \$4759 VGND sky130_fd_sc_hd__or2b_1
X$3324 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3331 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3332 VGND \$4761 \$4845 \$4406 \$4870 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3333 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3334 VGND \$4761 \$4821 \$4813 \$4871 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3336 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3337 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3340 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3341 VGND \$4761 \$4848 \$4813 \$4872 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3342 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3343 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3345 VPWR VGND \$4707 \$542 \$4857 \$4849 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3346 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3347 VPWR VGND VPWR \$4857 \$3122 VGND sky130_fd_sc_hd__inv_4
X$3348 VGND \$4353 \$4874 \$4850 \$4873 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3349 VPWR VGND VPWR \$4480 \$4874 VGND sky130_fd_sc_hd__inv_2
X$3350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3352 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3357 VGND \$4764 \$4839 \$4765 \$4875 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3358 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3361 VPWR VGND \$4899 \$184 \$4876 \$4888 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3362 VPWR VGND VPWR \$4173 \$4876 VGND sky130_fd_sc_hd__inv_2
X$3363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3365 VPWR \$4889 VGND \$1561 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$3366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3367 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3368 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3371 VGND \$4353 \$4840 \$4427 \$4858 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3374 VPWR \$2846 \$4877 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$3375 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3376 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3380 VGND \$2989 \$4830 \$4828 \$4859 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3382 VPWR \$4860 VGND VPWR \$4878 \$4492 \$3890 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$3383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3384 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3385 VPWR \$4831 VGND VPWR \$3036 VGND sky130_fd_sc_hd__clkbuf_1
X$3386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3387 VPWR VGND mgmt_gpio_oeb[14] VPWR \$4832 VGND sky130_fd_sc_hd__buf_2
X$3388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3391 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3393 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3395 VPWR \$481 \$810 \$439 VPWR VGND \$597 \$790 VGND sky130_fd_sc_hd__or4_1
X$3396 VGND \$733 \$781 \$801 \$748 \$598 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4bb_1
X$3397 VGND \$811 \$564 \$780 \$802 \$597 \$748 VPWR VPWR VGND
+ sky130_fd_sc_hd__a41o_1
X$3398 VGND \$802 \$739 \$790 \$439 \$599 VPWR VPWR VGND sky130_fd_sc_hd__o31a_1
X$3399 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3401 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3402 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3404 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3405 VPWR \$709 \$780 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3406 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3410 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3411 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3412 VPWR VGND VPWR \$812 \$227 VGND sky130_fd_sc_hd__inv_2
X$3413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3414 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3415 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3417 VPWR VGND \$701 \$200 \$791 \$814 \$711 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3419 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3420 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3421 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3422 VPWR VGND \$792 \$293 \$783 \$761 \$793 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3424 VPWR VGND \$792 \$294 \$794 \$817 \$793 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3425 VPWR VGND \$783 \$818 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$3426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3427 VPWR \$742 VGND \$1266 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$3428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3429 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3432 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3433 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3436 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3439 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3440 VGND \$516 \$860 \$605 \$797 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3442 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3443 VPWR VGND \$627 \$183 \$798 \$831 \$607 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3444 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3445 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3446 VPWR VGND VPWR \$796 \$737 VGND sky130_fd_sc_hd__inv_2
X$3447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3449 VGND \$516 \$772 \$771 \$786 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3450 VPWR \$773 VGND \$379 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$3451 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3452 VPWR VGND \$713 \$183 \$799 \$832 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3453 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3456 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3457 VGND \$516 \$849 \$435 \$805 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3458 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3459 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3460 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3461 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3462 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3463 VGND \$516 \$775 \$466 \$788 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3464 VGND \$516 \$823 \$466 \$806 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3465 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3466 VGND \$692 \$789 \$787 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3467 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3468 VGND \$824 \$562 \$930 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3470 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3471 VGND \$516 \$825 \$541 \$807 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3474 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3475 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3476 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3477 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3478 VPWR VGND VPWR \$776 \$808 VGND sky130_fd_sc_hd__inv_2
X$3479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3480 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3481 VPWR VGND \$826 VPWR mgmt_gpio_in[1] VGND sky130_fd_sc_hd__clkbuf_4
X$3482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3483 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3484 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3485 VPWR VGND VPWR \$840 \$827 VGND sky130_fd_sc_hd__inv_2
X$3486 VPWR \$827 VGND VPWR sram_ro_data[4] VGND sky130_fd_sc_hd__clkbuf_1
X$3487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3488 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3489 VPWR \$828 VGND VPWR \$810 VGND sky130_fd_sc_hd__clkbuf_1
X$3490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3491 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3492 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3495 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3496 VPWR \$813 VGND VPWR \$829 VGND sky130_fd_sc_hd__clkbuf_1
X$3497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3498 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3499 VGND \$655 \$854 \$237 \$841 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3500 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3502 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3503 VPWR VGND VPWR \$443 \$429 VGND sky130_fd_sc_hd__inv_2
X$3504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3506 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3507 VPWR VGND \$443 \$354 \$484 \$843 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3509 VPWR VGND \$429 VPWR \$845 VGND sky130_fd_sc_hd__clkbuf_4
X$3510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3511 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3512 VPWR \$845 VGND \$686 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$3513 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3515 VGND \$655 \$791 \$922 \$814 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3517 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3518 VPWR VGND VPWR \$792 \$793 VGND sky130_fd_sc_hd__inv_2
X$3519 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3520 VPWR \$846 VGND \$816 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$3521 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3522 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3523 VGND \$655 \$794 \$196 \$817 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3526 VPWR VGND \$794 \$815 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$3527 VGND \$820 \$337 \$818 \$816 \$325 \$782 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3529 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3530 VPWR VGND \$602 \$281 \$847 \$830 \$674 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3535 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3536 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3537 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3538 VGND \$516 \$798 \$771 \$831 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3542 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3545 VGND \$516 \$799 \$435 \$832 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3547 VPWR \$833 VGND \$848 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$3548 VPWR VGND \$714 VPWR \$833 VGND sky130_fd_sc_hd__clkbuf_4
X$3549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3550 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3551 VPWR VGND \$713 \$411 \$849 \$805 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3552 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3553 VGND \$834 \$849 \$821 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3554 VGND \$516 \$835 \$466 \$850 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3555 VGND \$822 \$835 \$834 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3557 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3558 VGND \$765 \$823 \$941 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3559 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3560 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3561 VGND \$766 \$289 \$789 \$824 \$851 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3563 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3564 VGND \$807 \$289 \$825 \$836 \$837 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3566 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3567 VGND \$707 \$825 \$838 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3568 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3569 VGND \$516 \$322 \$541 \$852 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$3570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3572 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3575 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3578 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3579 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3580 VPWR \$310 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3581 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3582 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3583 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3585 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3586 VPWR \$311 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3587 VPWR \$311 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3589 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3590 VPWR \$311 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3591 VPWR \$302 VGND \$311 \$308 VPWR VGND sky130_fd_sc_hd__or2_1
X$3592 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3593 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3594 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3595 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3596 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3599 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3601 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3603 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3604 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3605 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3606 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3608 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3610 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3611 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3613 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3618 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3619 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3622 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3623 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3625 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3627 VGND \$318 \$303 \$319 \$326 \$258 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3629 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3632 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3635 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3636 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3638 VGND \$321 \$189 \$433 \$320 \$185 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3639 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3642 VGND \$272 \$248 \$305 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3643 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3644 VGND \$206 \$290 \$246 \$298 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3645 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3646 VGND \$233 \$323 \$644 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3647 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3648 VGND \$250 \$289 \$222 \$324 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3650 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3651 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3652 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3654 VGND \$300 \$252 \$268 \$304 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$3655 VPWR VGND \$291 \$184 \$268 \$224 \$292 VPWR VGND sky130_fd_sc_hd__a22o_1
X$3656 VPWR \$291 \$292 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3658 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3659 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3660 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3662 VPWR VGND VPWR \$301 \$306 VGND sky130_fd_sc_hd__inv_2
X$3663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3667 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3668 VGND \$328 \$310 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$3669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3671 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3672 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3673 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3678 VPWR \$331 VGND VPWR \$329 VGND sky130_fd_sc_hd__clkbuf_1
X$3679 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3680 VGND \$329 \$194 \$183 \$273 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3681 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3682 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3683 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3684 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3686 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3687 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3688 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3690 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3691 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3694 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3695 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3696 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3697 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3698 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3699 VGND \$336 \$316 \$320 \$325 \$314 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3701 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3702 VPWR \$337 VGND VPWR \$312 \$353 \$285 \$326 VGND sky130_fd_sc_hd__o22a_1
X$3703 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3704 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3705 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3706 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3710 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3711 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3713 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3714 VPWR \$355 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3716 VPWR \$277 VGND \$319 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$3717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3720 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3726 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3727 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3728 VGND \$206 \$339 \$435 \$349 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3729 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3730 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3731 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3732 VGND \$327 \$290 \$330 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3733 VGND \$299 \$289 \$323 \$327 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$3734 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3736 VGND \$206 \$341 \$246 \$340 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3737 VGND \$324 \$341 \$502 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3740 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3741 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3744 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3746 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3749 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3751 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3752 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3754 VGND \$1667 \$1684 \$1376 \$1652 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$3755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3756 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3757 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3758 VPWR \$1642 \$1618 VGND VPWR VGND sky130_fd_sc_hd__clkdlybuf4s25_1
X$3759 VPWR VGND \$1514 \$1786 \$1633 \$1642 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3762 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3763 VGND \$1653 \$1580 \$1634 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3764 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3765 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3766 VPWR VGND VPWR \$1609 \$1620 VGND sky130_fd_sc_hd__inv_2
X$3767 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3768 VGND \$1525 \$1580 \$1620 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3769 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3770 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3772 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3779 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3780 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3781 VPWR \$1621 VGND \$1643 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$3782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3783 VGND \$856 \$1658 \$1370 \$1656 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3784 VGND \$856 \$1622 \$463 \$1638 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3785 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3786 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3787 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3788 VPWR \$1598 VGND VPWR \$1643 \$1425 VGND sky130_fd_sc_hd__or2_4
X$3789 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3791 VPWR \$1657 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3792 VGND \$1659 \$1600 \$1644 \$1198 \$1556 \$1655 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3793 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3794 VPWR \$1598 VGND VPWR \$1645 \$1420 VGND sky130_fd_sc_hd__or2_4
X$3795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3796 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3799 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3800 VGND \$1646 \$1615 \$1465 \$325 \$360 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$3801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3804 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3806 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3808 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3809 VPWR VGND \$1303 \$1179 \$1647 \$1660 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3811 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3812 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3813 VPWR VGND \$1303 \$184 \$1648 \$1661 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3817 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3819 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3820 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3821 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3822 VGND \$1152 \$1649 \$541 \$1629 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3823 VGND \$1630 \$895 \$1308 \$1662 \$1649 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$3824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3825 VPWR \$1663 VPWR VGND \$1308 \$1650 VGND sky130_fd_sc_hd__or2_2
X$3826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3828 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3829 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3831 VGND \$516 \$1664 \$1273 \$1641 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3832 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3833 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3834 VPWR VGND \$1311 \$411 \$1651 \$1665 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3835 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3837 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3839 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3841 VPWR \$1682 VGND VPWR sram_ro_data[19] VGND sky130_fd_sc_hd__clkbuf_1
X$3842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3843 VPWR \$1667 VGND VPWR \$1632 VGND sky130_fd_sc_hd__clkbuf_1
X$3844 VPWR VGND \$1514 \$1683 \$1684 \$1652 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3845 VGND \$1683 \$907 \$1498 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3846 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3847 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3848 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3849 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3851 VPWR \$1685 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$3852 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3853 VPWR VGND \$1053 \$1653 \$1620 \$1686 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3855 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3856 VPWR VGND \$1053 \$1687 \$1487 \$1688 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3858 VPWR \$1689 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$3859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3860 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3861 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3863 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3866 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3867 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3870 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3871 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3872 VGND \$1668 \$1059 \$1034 \$1654 \$1643 \$1443 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$3873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3875 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3876 VPWR VGND \$1567 \$294 \$1658 \$1656 \$1568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3877 VPWR VGND VPWR \$1675 \$1658 VGND sky130_fd_sc_hd__inv_2
X$3878 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3879 VPWR \$1690 VGND VPWR \$1675 \$1613 \$274 \$325 VGND
+ sky130_fd_sc_hd__o22a_1
X$3880 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3882 VPWR VGND VPWR \$1639 \$1622 VGND sky130_fd_sc_hd__inv_2
X$3883 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3884 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3886 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3887 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3888 VPWR VGND VPWR \$1670 \$1657 \$1659 \$820 \$1669 VGND
+ sky130_fd_sc_hd__and4_1
X$3889 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3890 VPWR \$1692 VGND \$1034 \$1434 VPWR VGND sky130_fd_sc_hd__or2_1
X$3891 VPWR \$1490 VGND VPWR \$1676 \$1264 VGND sky130_fd_sc_hd__or2_4
X$3892 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3893 VPWR \$1677 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3894 VPWR \$1693 VGND VPWR \$784 \$744 \$1677 \$1588 VGND
+ sky130_fd_sc_hd__o22a_1
X$3895 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3896 VPWR \$1694 VGND VPWR \$1163 \$1271 \$1678 \$1300 VGND
+ sky130_fd_sc_hd__o22a_1
X$3897 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3898 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3900 VPWR \$1615 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$3901 VPWR \$1696 VGND VPWR \$1121 \$1562 \$1639 \$1613 VGND
+ sky130_fd_sc_hd__o22a_1
X$3902 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3903 VGND \$1718 \$589 \$265 \$433 \$1645 \$1616 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3904 VPWR VGND VPWR \$1699 \$1698 \$1697 \$940 \$1082 VGND
+ sky130_fd_sc_hd__and4_1
X$3905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3908 VPWR VGND VPWR \$1778 \$1626 VGND sky130_fd_sc_hd__inv_2
X$3909 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3911 VGND \$1152 \$1647 \$1627 \$1660 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$3912 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3913 VGND \$1152 \$1648 \$1203 \$1661 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3915 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3916 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3917 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3918 VPWR VGND VPWR \$1702 \$1593 VGND sky130_fd_sc_hd__inv_2
X$3919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3920 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3921 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3922 VPWR \$1672 VPWR VGND \$1322 \$1128 \$1679 VGND sky130_fd_sc_hd__or3_1
X$3923 VGND \$1672 \$2670 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$3924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3925 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3926 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3927 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3928 VPWR \$1798 VPWR VGND \$1531 \$1574 \$1673 VGND sky130_fd_sc_hd__or3_2
X$3929 VPWR VGND VPWR \$1673 \$1649 VGND sky130_fd_sc_hd__inv_2
X$3930 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3931 VGND \$1706 \$1663 \$895 \$1650 \$1797 \$672 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$3932 VPWR \$1798 VPWR VGND \$1346 \$1650 VGND sky130_fd_sc_hd__or2_2
X$3933 VPWR VGND VPWR \$1650 \$1662 VGND sky130_fd_sc_hd__inv_2
X$3934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3935 VPWR VGND \$1680 \$411 \$1707 \$1708 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3937 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3938 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3940 VPWR VGND VPWR \$1664 \$1225 VGND sky130_fd_sc_hd__inv_4
X$3941 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3942 VGND \$516 \$1651 \$1273 \$1665 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3943 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3944 VGND \$1710 \$1594 \$1595 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$3945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3946 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3947 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3948 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3950 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3951 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3952 VPWR \$2833 VGND \$2424 VPWR \$1979 VGND sky130_fd_sc_hd__nor2_1
X$3953 VPWR \$2834 VGND \$2320 VPWR \$2537 VGND sky130_fd_sc_hd__nor2_1
X$3954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3955 VPWR \$2712 VPWR VGND \$2835 \$2834 \$2676 VGND sky130_fd_sc_hd__or3_1
X$3956 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3957 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3958 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3961 VPWR \$2816 VGND \$2659 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$3962 VPWR \$2817 VPWR VGND \$2168 \$2816 VGND sky130_fd_sc_hd__nand2_1
X$3963 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3966 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3967 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3968 VPWR VGND VPWR \$2836 \$2744 VGND sky130_fd_sc_hd__inv_2
X$3969 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3971 VPWR \$2837 VGND \$2745 \$2259 VPWR VGND sky130_fd_sc_hd__or2_1
X$3972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3975 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3976 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3977 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3978 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$3979 VPWR \$2719 \$2732 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$3980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$3981 VGND \$856 \$2839 \$2556 \$2838 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$3982 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3983 VPWR VGND VPWR \$2818 \$2733 VGND sky130_fd_sc_hd__inv_2
X$3984 VPWR VGND VPWR \$2747 \$2839 VGND sky130_fd_sc_hd__inv_2
X$3985 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$3986 VPWR VGND \$2703 \$183 \$2764 \$2799 \$2705 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$3987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$3989 VGND \$2820 \$2800 \$2819 \$2358 \$2274 \$2840 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3991 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$3992 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$3993 VGND \$2821 \$2820 \$495 \$785 \$2220 \$2747 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3994 VGND \$2822 \$2802 \$2821 VPWR \$609 VPWR VGND sky130_fd_sc_hd__nand3_4
X$3995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$3996 VGND \$2823 \$2527 \$2684 \$2043 \$1914 \$762 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$3997 VGND \$1123 \$2818 \$2778 \$2386 \$2841 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$3998 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$3999 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4000 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4002 VPWR \$1264 VGND VPWR \$2614 \$1571 VGND sky130_fd_sc_hd__or2_4
X$4003 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4005 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4006 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4007 VPWR \$2824 VGND VPWR \$1294 \$1776 \$3444 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$4008 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4009 VGND \$2825 \$2824 \$2752 \$1715 \$1754 \$1330 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4010 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4011 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4012 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4013 VGND \$2827 \$2826 \$2561 \$2116 \$1536 \$1481 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4014 VPWR VGND VPWR \$2844 \$2825 \$2827 \$2828 \$2842 VGND
+ sky130_fd_sc_hd__and4_1
X$4015 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4016 VPWR \$2843 VGND VPWR \$2502 \$2254 \$2669 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$4017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4018 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4019 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4022 VGND \$2810 \$2845 \$1373 \$2525 \$2458 \$2829 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4023 VPWR \$2845 VGND VPWR \$1855 \$2456 \$2846 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$4024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4025 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4026 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4027 VPWR \$2847 VGND VPWR \$500 \$2045 \$2671 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$4028 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4029 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4031 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4032 VPWR \$2831 VGND \$2785 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$4033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4034 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4036 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4037 VPWR VGND \$2832 \$1880 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4039 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4040 VPWR VGND \$2711 VPWR \$2831 VGND sky130_fd_sc_hd__clkbuf_4
X$4041 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4043 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4047 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4048 VPWR \$2849 VGND VPWR \$2856 VGND sky130_fd_sc_hd__clkbuf_1
X$4049 VPWR VGND mgmt_gpio_oeb[7] VPWR \$2849 VGND sky130_fd_sc_hd__buf_2
X$4050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4051 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4052 VGND trap \$2869 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$4053 VPWR \$2857 \$2622 \$2890 VPWR VGND \$2833 \$2834 VGND
+ sky130_fd_sc_hd__or4_1
X$4054 VPWR \$2676 VGND \$2833 \$2870 VPWR VGND sky130_fd_sc_hd__or2_1
X$4055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4057 VPWR \$2858 VGND \$2659 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$4058 VGND \$2740 \$2816 \$2858 \$2871 \$2891 \$2741 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$4059 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4060 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4062 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4063 VPWR \$2661 VGND \$2514 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$4064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4065 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4066 VPWR \$2874 VGND \$2836 \$2017 VPWR VGND sky130_fd_sc_hd__or2_1
X$4067 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4069 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4071 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4072 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4073 VPWR VGND \$2775 \$183 \$2875 \$2851 \$2776 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4076 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4077 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4079 VPWR VGND VPWR \$1325 \$2859 VGND sky130_fd_sc_hd__inv_2
X$4080 VPWR VGND \$2876 \$294 \$2839 \$2838 \$2934 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4081 VPWR VGND VPWR \$2779 \$2778 VGND sky130_fd_sc_hd__inv_2
X$4082 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4083 VPWR VGND VPWR \$2749 \$2877 VGND sky130_fd_sc_hd__inv_2
X$4084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4086 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4087 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4088 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4090 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4092 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4093 VPWR \$2778 VPWR VGND \$1034 \$1445 VGND sky130_fd_sc_hd__or2_2
X$4094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4095 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4096 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4097 VPWR VGND VPWR \$2822 \$1764 \$2860 \$2823 \$2878 VGND
+ sky130_fd_sc_hd__and4_1
X$4098 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4099 VGND \$2852 \$2861 \$2840 \$2544 \$2545 \$2684 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4103 VPWR \$2788 VGND VPWR \$2781 \$2384 \$2806 \$1645 VGND
+ sky130_fd_sc_hd__o22a_1
X$4104 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4105 VPWR \$1329 VGND VPWR \$2789 \$1571 VGND sky130_fd_sc_hd__or2_4
X$4106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4107 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4108 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4109 VPWR \$2881 VGND VPWR \$1330 \$2724 \$2615 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$4110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4111 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4113 VPWR \$2826 VGND \$2007 \$2900 VPWR VGND sky130_fd_sc_hd__or2_1
X$4114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4115 VGND \$2842 \$2843 \$2806 \$2809 \$3218 \$2853 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4117 VPWR \$2882 VGND VPWR \$1023 \$2724 \$2854 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$4118 VGND \$2793 \$2882 \$1949 \$2369 \$2357 \$2862 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4120 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4121 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4123 VPWR \$2794 VGND VPWR \$2863 \$2544 \$2908 \$2545 VGND
+ sky130_fd_sc_hd__o22a_1
X$4124 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4125 VGND \$2755 \$1803 \$2005 \$2864 \$2865 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$4126 VPWR \$2864 VGND VPWR \$2866 \$2670 \$1221 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$4127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4128 VGND \$2884 \$2847 \$2923 \$2073 \$2096 \$2846 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4131 VGND \$2885 \$2867 \$1892 \$2809 \$3218 \$2829 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4133 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4135 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4136 VPWR VGND \$2633 \$1171 \$2868 \$2886 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4138 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4139 VPWR VGND \$2633 \$542 \$2855 \$2887 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4140 VGND \$1152 \$2855 \$2450 \$2887 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$4141 VPWR VGND \$2694 \$411 \$2832 \$2888 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4142 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4143 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4146 VGND \$1152 \$2963 \$2232 \$2889 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4150 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4151 VPWR \$2856 VGND VPWR \$2906 VGND sky130_fd_sc_hd__clkbuf_1
X$4152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4156 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4157 VPWR \$5456 VGND VPWR \$5189 \$5439 \$5448 \$1829 VGND
+ sky130_fd_sc_hd__o22a_1
X$4158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4160 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4162 VPWR VGND \$5448 VPWR \$5363 VGND sky130_fd_sc_hd__clkbuf_4
X$4163 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4166 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4168 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4169 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4170 VPWR \$5440 VGND \$4474 VPWR \$5449 VGND sky130_fd_sc_hd__nor2_1
X$4171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4175 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4176 VGND \$5442 \$5450 \$4106 \$5441 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4177 VGND \$5443 \$5486 \$4106 \$5459 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4180 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4186 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4187 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4189 VPWR VGND \$5097 \$3694 \$5436 \$5460 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4190 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4191 VGND \$2777 \$5462 \$5408 \$5451 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4192 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4194 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4195 VPWR VGND \$5461 \$3236 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4197 VGND \$4761 \$5437 \$4994 \$5444 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4200 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4201 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4203 VPWR VGND VPWR \$3936 \$5452 VGND sky130_fd_sc_hd__inv_2
X$4204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4207 VPWR \$4560 \$5453 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4208 VPWR VGND \$5332 \$4774 \$5453 \$5478 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4209 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4212 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4213 VPWR VGND \$5463 VPWR \$5263 VGND sky130_fd_sc_hd__clkbuf_4
X$4214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4217 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4218 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4219 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4220 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4222 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4223 VPWR \$5344 \$5312 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4226 VPWR \$2863 \$5490 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$4227 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4228 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4230 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4231 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4232 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4233 VGND \$4764 \$5464 \$5298 \$5445 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4235 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4236 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4237 VPWR \$5438 VGND VPWR \$5429 \$4724 \$5454 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$4238 VGND \$5454 \$1892 mgmt_gpio_out[17] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$4239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4241 VGND \$5189 \$5002 \$5456 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$4242 VPWR \$5492 VGND VPWR \$5145 \$5439 \$5448 \$907 VGND
+ sky130_fd_sc_hd__o22a_1
X$4243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4245 VPWR \$5466 \$5457 VGND \$5502 VPWR \$4833 VGND sky130_fd_sc_hd__nor3_1
X$4246 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4247 VPWR \$5415 VPWR VGND \$5466 \$5482 \$5467 VGND sky130_fd_sc_hd__or3_1
X$4248 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4249 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4251 VPWR VPWR VGND \$4892 \$5468 \$4733 \$5406 VGND sky130_fd_sc_hd__a21bo_2
X$4252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4253 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4254 VPWR \$5483 VGND VPWR \$4576 \$5469 VGND sky130_fd_sc_hd__or2_4
X$4255 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4256 VPWR \$5470 VPWR VGND \$5326 \$5471 \$5458 VGND sky130_fd_sc_hd__or3_2
X$4257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4258 VPWR VGND VPWR \$5220 \$5467 VGND sky130_fd_sc_hd__inv_2
X$4259 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4260 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4261 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4262 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4265 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4267 VPWR VGND \$5504 \$5485 \$5486 \$5459 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4268 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4269 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4270 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4277 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4280 VPWR VGND \$5192 \$411 \$5473 \$5472 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4282 VPWR VGND \$5473 \$3714 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4283 VGND \$4374 \$5165 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$4284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4285 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4286 VPWR VGND \$5097 \$1594 \$5461 \$5474 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4287 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4288 VGND \$2777 \$5461 \$5408 \$5474 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4291 VPWR VGND VPWR \$3436 \$5475 VGND sky130_fd_sc_hd__inv_2
X$4292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4294 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4297 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4298 VGND \$4761 \$5452 \$5367 \$5476 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4299 VPWR VGND \$5477 \$2666 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4300 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4301 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4302 VGND \$4761 \$5453 \$5367 \$5478 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4305 VPWR VGND VPWR \$3771 \$5499 VGND sky130_fd_sc_hd__inv_2
X$4306 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4308 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4309 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4310 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4311 VPWR VGND VPWR \$5332 \$5391 VGND sky130_fd_sc_hd__inv_2
X$4312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4313 VPWR VGND \$5332 \$3694 \$5488 \$5487 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4316 VPWR VGND VPWR \$3543 \$5479 VGND sky130_fd_sc_hd__inv_2
X$4317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4318 VPWR VGND \$5344 \$411 \$5479 \$5489 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4321 VPWR VGND VPWR \$5480 \$2691 VGND sky130_fd_sc_hd__inv_4
X$4322 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4323 VPWR VGND \$5344 \$3694 \$5490 \$5481 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4324 VGND \$4764 \$5490 \$5334 \$5481 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$4325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4328 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4329 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4330 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4331 VPWR VGND \$5335 \$1594 \$5464 \$5445 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4335 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4336 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4337 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4338 VPWR \$5491 VGND VPWR \$5446 VGND sky130_fd_sc_hd__clkbuf_1
X$4339 VPWR VGND mgmt_gpio_oeb[17] VPWR \$5491 VGND sky130_fd_sc_hd__buf_2
X$4340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4341 VPWR \$2012 VGND VPWR sram_ro_data[24] VGND sky130_fd_sc_hd__clkbuf_1
X$4342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4343 VPWR \$2038 VGND VPWR sram_ro_data[25] VGND sky130_fd_sc_hd__clkbuf_1
X$4344 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4346 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4347 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4351 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4353 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4354 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4358 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4359 VPWR VGND \$1725 \$2070 \$2082 \$2092 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4361 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4363 VPWR VGND \$1923 \$183 \$2083 \$2093 \$1924 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4367 VPWR VGND \$1752 \$294 \$2084 \$2094 \$1774 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4368 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4369 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4370 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4371 VGND \$856 \$2071 \$1861 \$2085 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4372 VGND \$856 \$2095 \$1863 \$2086 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4374 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4376 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4377 VGND \$2074 \$2087 \$702 \$2073 \$2096 \$2072 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4378 VPWR \$1490 VGND VPWR \$2031 \$1420 VGND sky130_fd_sc_hd__or2_4
X$4379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4380 VGND \$2097 \$2075 \$2088 \$2043 \$1914 \$726 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4381 VPWR \$2075 VGND VPWR \$2076 \$1966 \$1691 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$4382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4383 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4384 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4387 VGND \$2227 \$703 \$2045 \$1955 \$1529 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$4388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4389 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4390 VGND \$2077 \$882 \$2005 \$2098 \$2032 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$4391 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4393 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4394 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4396 VGND \$2021 \$2066 \$2047 \$2048 \$646 \$2099 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$4397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4400 VGND \$2100 \$1990 \$2089 \$2031 \$2113 \$2066 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4403 VPWR VGND VPWR \$2049 \$2050 VGND sky130_fd_sc_hd__inv_2
X$4404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4405 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4406 VGND \$1152 \$2051 \$1203 \$2067 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4409 VPWR \$2079 VPWR VGND \$1438 \$1882 \$1705 VGND sky130_fd_sc_hd__or3_1
X$4410 VGND \$2052 \$2135 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$4411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4412 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4413 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4414 VPWR \$1971 VGND \$2080 \$1782 VPWR VGND sky130_fd_sc_hd__or2_1
X$4415 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4416 VGND \$2081 \$1065 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$4417 VGND \$1994 \$3218 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$4418 VPWR \$2054 VGND \$1801 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$4419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4420 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4421 VGND \$1152 \$2101 \$1273 \$2090 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4425 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4426 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4430 VPWR \$2102 VGND VPWR \$2033 VGND sky130_fd_sc_hd__clkbuf_1
X$4431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4432 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4435 VPWR \$2129 VGND VPWR sram_ro_data[26] VGND sky130_fd_sc_hd__clkbuf_1
X$4436 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4439 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4440 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4441 VPWR \$2130 VGND \$1960 \$1979 VPWR VGND sky130_fd_sc_hd__or2_1
X$4442 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4443 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4444 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4445 VPWR \$2131 VGND \$2119 VPWR \$1999 VGND sky130_fd_sc_hd__nor2_1
X$4446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4448 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4449 VPWR \$2133 VGND \$1981 \$2017 VPWR VGND sky130_fd_sc_hd__or2_1
X$4450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4451 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4452 VPWR \$2104 VGND \$2026 VPWR \$1998 VGND sky130_fd_sc_hd__nor2_1
X$4453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4454 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4455 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4456 VGND \$856 \$2083 \$1750 \$2093 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4458 VPWR VGND \$1923 \$293 \$2134 \$2157 \$1924 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4459 VPWR \$2121 \$2083 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4460 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4462 VPWR \$1744 \$2134 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4464 VGND \$856 \$2084 \$1861 \$2094 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4465 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4466 VPWR VGND \$2120 \$200 \$2071 \$2085 \$2106 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4468 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4469 VPWR VGND \$2120 \$183 \$2095 \$2086 \$2106 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4470 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4471 VPWR VGND VPWR \$2076 \$2095 VGND sky130_fd_sc_hd__inv_2
X$4472 VPWR \$2218 VGND VPWR \$1265 \$2135 \$1852 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$4473 VPWR \$2108 VGND VPWR \$1192 \$2135 \$2121 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$4474 VGND \$2136 \$2108 \$2122 \$1065 \$880 \$2123 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4476 VGND \$2124 \$2137 \$2125 VPWR \$570 VPWR VGND sky130_fd_sc_hd__nand3_4
X$4477 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4479 VPWR \$2109 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$4480 VPWR VGND VPWR \$2124 \$1866 \$2138 \$2097 \$2109 VGND
+ sky130_fd_sc_hd__and4_1
X$4481 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4482 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4483 VPWR \$2139 VGND VPWR \$2121 \$1967 \$1691 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$4484 VGND \$2140 \$2139 \$784 \$1953 \$1987 \$1024 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4486 VPWR \$2110 VGND VPWR \$1948 \$1713 \$1023 \$859 VGND
+ sky130_fd_sc_hd__o22a_1
X$4487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4488 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4489 VGND \$1790 \$2110 \$2018 \$1729 \$1625 \$2111 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4492 VPWR \$2112 VGND VPWR \$1024 \$1956 \$1820 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$4493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4494 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4495 VPWR \$2141 VGND VPWR \$1628 \$1198 \$1611 \$1643 VGND
+ sky130_fd_sc_hd__o22a_1
X$4496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4497 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4498 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4499 VGND \$869 \$2100 \$2114 \$2142 \$1876 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$4500 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4501 VPWR VGND \$2049 \$183 \$2143 \$2144 \$2050 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4503 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4504 VPWR \$1335 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$4505 VPWR \$2115 \$1333 VPWR \$2020 VGND \$2113 \$1335 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$4506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4507 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4508 VPWR VGND VPWR \$2145 \$3218 \$1957 \$2073 \$2116 VGND
+ sky130_fd_sc_hd__and4_1
X$4509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4510 VPWR VGND VPWR \$1136 \$2146 \$2145 \$844 \$1766 VGND
+ sky130_fd_sc_hd__and4_1
X$4511 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4513 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4514 VPWR \$2147 VPWR VGND \$1814 \$1663 \$1766 VGND sky130_fd_sc_hd__or3_1
X$4515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4516 VPWR \$2148 VGND \$1813 \$1782 VPWR VGND sky130_fd_sc_hd__or2_1
X$4517 VGND \$2126 \$844 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$4518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4519 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4520 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4521 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4522 VPWR \$2149 \$1183 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4523 VGND \$2149 \$1406 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$4524 VPWR VGND \$1680 \$1179 \$2101 \$2090 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4527 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4528 VPWR \$1083 VGND VPWR \$2117 \$2149 VGND sky130_fd_sc_hd__or2_4
X$4529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4530 VPWR VGND \$2127 \$411 \$2151 \$2185 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4535 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4536 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4537 VPWR \$2152 VGND VPWR \$2102 VGND sky130_fd_sc_hd__clkbuf_1
X$4538 VPWR VGND mgmt_gpio_oeb[5] VPWR \$2152 VGND sky130_fd_sc_hd__buf_2
X$4539 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4540 VPWR \$853 VGND VPWR sram_ro_data[5] VGND sky130_fd_sc_hd__clkbuf_1
X$4541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4542 VPWR \$875 VGND VPWR \$863 VGND sky130_fd_sc_hd__clkbuf_1
X$4543 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4544 VPWR \$863 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$4545 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4547 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4548 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4549 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4550 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4552 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4553 VPWR \$865 VPWR VGND \$854 \$599 \$235 VGND sky130_fd_sc_hd__or3_1
X$4554 VPWR \$878 VGND VPWR \$898 VGND sky130_fd_sc_hd__clkbuf_1
X$4555 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4556 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4557 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4559 VPWR \$829 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$4560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4561 VPWR \$841 VGND VPWR \$866 VGND sky130_fd_sc_hd__clkbuf_1
X$4562 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4563 VGND \$866 \$854 \$183 \$867 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4566 VPWR VGND \$443 \$281 \$343 \$855 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4567 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4568 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4569 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4570 VPWR VGND \$443 \$411 \$461 \$879 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4572 VGND \$856 \$484 \$239 \$843 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$4573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4575 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4576 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4578 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4579 VPWR VGND \$791 \$868 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4580 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4581 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4582 VPWR VPWR VGND \$846 \$793 VGND sky130_fd_sc_hd__clkbuf_2
X$4583 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4585 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4586 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4587 VGND \$655 \$858 \$196 \$857 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4589 VGND \$655 \$847 \$961 \$830 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4590 VPWR VGND \$847 \$882 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4592 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4594 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4595 VPWR \$885 VGND \$859 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$4596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4597 VPWR VGND \$912 \$200 \$860 \$797 \$893 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4600 VPWR VGND \$860 \$803 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$4601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4602 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4603 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4604 VPWR VGND VPWR \$819 \$798 VGND sky130_fd_sc_hd__inv_2
X$4605 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4606 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4607 VGND \$869 \$287 \$803 \$859 \$433 \$249 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4609 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4610 VPWR VGND VPWR \$861 \$772 VGND sky130_fd_sc_hd__inv_2
X$4611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4612 VPWR VGND VPWR \$870 \$799 VGND sky130_fd_sc_hd__inv_2
X$4613 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4614 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4615 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4616 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4617 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4618 VPWR VGND VPWR \$871 \$849 VGND sky130_fd_sc_hd__inv_2
X$4619 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4620 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4621 VPWR \$862 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$4622 VGND \$787 \$849 \$862 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4624 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4625 VGND \$850 \$289 \$835 \$887 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$4626 VGND \$887 \$775 \$872 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4628 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4629 VGND \$806 \$289 \$823 \$888 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$4630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4633 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4634 VPWR VGND VPWR \$289 \$851 VGND sky130_fd_sc_hd__inv_4
X$4635 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4637 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4638 VPWR VGND VPWR \$289 \$837 VGND sky130_fd_sc_hd__inv_4
X$4639 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4642 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4646 VPWR VGND mgmt_gpio_oeb[1] VPWR \$873 VGND sky130_fd_sc_hd__buf_2
X$4647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4649 VGND \$875 \$906 \$381 \$896 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4651 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4652 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4653 VPWR \$876 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$4654 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4655 VPWR \$877 VGND VPWR \$876 VGND sky130_fd_sc_hd__clkbuf_1
X$4656 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4657 VGND \$878 \$1015 \$387 \$751 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$4658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4661 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4663 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4664 VGND \$856 \$343 \$891 \$855 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$4665 VGND \$856 \$461 \$891 \$879 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$4666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4667 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4671 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4673 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4674 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4678 VPWR VGND \$892 \$293 \$858 \$857 \$911 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4681 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4682 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4684 VGND \$655 \$884 \$605 \$883 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4685 VPWR VGND \$912 \$184 \$884 \$883 \$893 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4686 VPWR VGND \$893 VPWR \$885 VGND sky130_fd_sc_hd__clkbuf_4
X$4687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4688 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4689 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4690 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4693 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4694 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4696 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4697 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4698 VGND \$886 \$730 \$929 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4699 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4700 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4701 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4702 VPWR VGND \$713 \$294 \$894 \$901 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$4703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4704 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4705 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4706 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4711 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4712 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4714 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4718 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4720 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4723 VPWR \$889 VPWR VGND \$902 \$808 VGND sky130_fd_sc_hd__or2_2
X$4724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4726 VPWR VGND VPWR \$904 \$759 VGND sky130_fd_sc_hd__inv_2
X$4727 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4728 VPWR \$904 \$903 \$915 VPWR VGND \$997 \$698 VGND sky130_fd_sc_hd__or4_1
X$4729 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4730 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4731 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4732 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4733 VPWR VGND VPWR \$1312 \$1111 VGND sky130_fd_sc_hd__inv_2
X$4734 VGND \$1313 \$1292 \$381 \$1277 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4736 VGND \$1269 \$1292 \$780 \$828 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4738 VGND \$1280 \$564 \$381 \$1254 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_4
X$4739 VPWR \$1270 VGND VPWR \$565 VGND sky130_fd_sc_hd__clkbuf_1
X$4740 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4741 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4742 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4744 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4745 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4749 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4752 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4753 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4754 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4755 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4756 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4757 VPWR \$1298 VGND VPWR \$1267 \$1297 \$958 \$1058 VGND
+ sky130_fd_sc_hd__o22a_1
X$4758 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4759 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4762 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4766 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4767 VPWR \$1264 VGND VPWR \$755 \$1034 VGND sky130_fd_sc_hd__or2_4
X$4768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4769 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4770 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4771 VPWR VGND \$912 \$411 \$1293 \$1285 \$893 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4773 VPWR VGND \$912 \$294 \$1250 \$1249 \$893 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4778 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4779 VGND \$1301 \$1124 \$1294 \$1300 \$379 \$861 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4782 VPWR \$1284 \$1252 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4784 VGND \$1152 \$1344 \$1203 \$1302 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4785 VPWR VGND \$1303 \$294 \$1287 \$1286 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4786 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4787 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4788 VGND \$1152 \$1305 \$1203 \$1304 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4789 VPWR \$1320 \$1305 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$4790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4791 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4792 VPWR VGND \$1170 \$184 \$1296 \$1321 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4794 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4795 VPWR VGND VPWR \$1306 \$1296 VGND sky130_fd_sc_hd__inv_2
X$4796 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4798 VPWR \$1260 VGND VPWR \$1882 \$1138 VGND sky130_fd_sc_hd__or2_4
X$4799 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4801 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4802 VGND \$516 \$1308 \$541 \$1307 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_2
X$4803 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4804 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4805 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4806 VGND \$516 \$1140 \$541 \$1309 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4808 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4809 VPWR VGND \$1311 \$1179 \$1289 \$1288 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4810 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4811 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4813 VPWR VGND \$1311 \$386 \$1275 \$1290 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4815 VGND \$516 \$1261 \$1274 \$1291 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4816 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4818 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4819 VPWR VGND VPWR \$1349 \$1276 VGND sky130_fd_sc_hd__inv_2
X$4820 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4821 VPWR \$1313 VGND VPWR \$1278 VGND sky130_fd_sc_hd__clkbuf_1
X$4822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4825 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4826 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4828 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4829 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4830 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4831 VPWR VGND \$1053 \$1336 \$1337 \$1314 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4832 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4833 VPWR VGND \$1145 VPWR \$1162 \$1351 \$1337 VGND sky130_fd_sc_hd__a21oi_1
X$4834 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4835 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4836 VPWR \$1338 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$4837 VPWR \$1352 VGND VPWR \$1338 VGND sky130_fd_sc_hd__clkbuf_1
X$4838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4839 VGND \$1369 \$1191 \$1324 \$1317 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$4840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4842 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4843 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4845 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4846 VPWR \$1339 VGND VPWR \$1312 \$1297 \$1831 \$923 VGND
+ sky130_fd_sc_hd__o22a_1
X$4847 VGND \$1316 \$1339 \$1325 \$1340 \$456 \$333 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4850 VGND \$1341 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__inv_8
X$4851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4852 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4853 VGND \$1327 \$1298 \$1282 \$1271 \$816 \$1004 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4854 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4855 VGND \$1353 \$1258 \$1317 \$1318 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$4856 VPWR \$1257 VGND VPWR \$1266 \$1342 VGND sky130_fd_sc_hd__or2_4
X$4857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4858 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4859 VGND \$1318 \$1329 \$1379 \$1353 \$1328 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$4860 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4861 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4862 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4863 VPWR \$1283 VGND VPWR \$1297 \$1248 VGND sky130_fd_sc_hd__or2_4
X$4864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4866 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4868 VPWR VGND \$912 \$354 \$1357 \$1319 \$893 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4870 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4871 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4872 VPWR \$1330 \$1250 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4874 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4875 VGND \$1152 \$1332 \$771 \$1343 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4876 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4877 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4879 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4880 VPWR VGND \$1303 \$183 \$1344 \$1302 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4882 VPWR VGND VPWR \$1294 \$1287 VGND sky130_fd_sc_hd__inv_2
X$4883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4884 VPWR VGND VPWR \$1303 \$1295 VGND sky130_fd_sc_hd__inv_2
X$4885 VPWR \$1359 VGND \$1300 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$4886 VPWR VGND \$1303 \$281 \$1305 \$1304 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4887 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4888 VPWR \$1331 VGND VPWR \$563 \$755 \$1320 \$1300 VGND
+ sky130_fd_sc_hd__o22a_1
X$4889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4890 VPWR \$1334 VGND VPWR \$1306 \$1198 \$255 \$755 VGND
+ sky130_fd_sc_hd__o22a_1
X$4891 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4894 VGND \$516 \$1296 \$993 \$1321 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4896 VPWR \$1260 VGND VPWR \$1360 \$1345 VGND sky130_fd_sc_hd__or2_4
X$4897 VPWR \$1137 VGND VPWR \$1322 \$1138 VGND sky130_fd_sc_hd__or2_4
X$4898 VPWR \$1322 \$1222 VGND \$1128 VPWR \$1011 VGND sky130_fd_sc_hd__nor3_1
X$4899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4901 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4902 VGND \$516 \$1374 \$541 \$1362 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$4903 VPWR \$1307 VGND VPWR \$1346 \$1011 \$1308 \$1323 VGND
+ sky130_fd_sc_hd__o22a_1
X$4904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4906 VPWR \$1323 VGND \$895 \$1140 VPWR VGND sky130_fd_sc_hd__or2_1
X$4907 VPWR \$672 \$1323 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4909 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4911 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4912 VGND \$1364 \$1179 \$1289 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$4913 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4914 VPWR VGND VPWR \$1311 \$1310 VGND sky130_fd_sc_hd__inv_2
X$4915 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4916 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4917 VGND mgmt_gpio_in[3] \$1333 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$4918 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4921 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4923 VPWR \$1505 \$1711 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4924 VPWR \$1722 \$1682 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4926 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4927 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4928 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4929 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4930 VPWR \$1723 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$4931 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4932 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4933 VGND \$1740 \$1620 \$1376 \$1686 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4935 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4936 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4938 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4939 VGND \$1742 \$1487 \$1376 \$1688 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$4940 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4941 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4942 VPWR VGND \$1725 \$1636 \$1741 \$1635 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4943 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4944 VPWR VGND \$1725 \$1324 \$1724 \$1674 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$4945 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4946 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4947 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4950 VPWR \$1726 VGND \$923 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$4951 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4952 VGND \$856 \$1728 \$1370 \$1727 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$4953 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4955 VPWR \$1691 \$1728 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$4956 VPWR \$1598 VGND VPWR \$1729 \$1059 VGND sky130_fd_sc_hd__or2_4
X$4957 VPWR \$1598 VGND VPWR \$1713 \$1444 VGND sky130_fd_sc_hd__or2_4
X$4958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4960 VGND \$1731 \$1690 \$1637 \$1643 \$1271 \$1256 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4961 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4962 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4963 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4964 VPWR \$1714 VGND VPWR \$1419 \$1776 \$818 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$4965 VGND \$1716 \$1714 \$1639 \$1715 \$1754 \$924 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4966 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4967 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4968 VPWR \$1671 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$4969 VGND \$1237 \$1668 \$1671 \$1645 \$1713 \$1691 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4971 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4972 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4973 VGND \$1732 \$1692 \$1730 \$1676 \$1554 \$1513 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4974 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4975 VGND \$1697 \$1744 \$1729 \$1694 \$1695 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$4976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$4977 VPWR \$1717 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$4978 VGND \$1695 \$581 \$1950 \$1340 \$1465 \$1717 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$4979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4980 VPWR VGND VPWR \$1719 \$1670 \$1733 \$1718 \$1734 VGND
+ sky130_fd_sc_hd__and4_1
X$4981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4982 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4983 VGND \$1703 \$1699 \$1719 VPWR \$907 VPWR VGND sky130_fd_sc_hd__nand3_4
X$4984 VGND \$1700 \$688 \$347 \$1692 \$1763 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$4985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4986 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4987 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$4988 VPWR VGND VPWR \$1678 \$1647 VGND sky130_fd_sc_hd__inv_2
X$4989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$4990 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4991 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$4992 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$4993 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$4994 VPWR VGND VPWR \$1720 \$1648 VGND sky130_fd_sc_hd__inv_2
X$4995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$4996 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$4997 VGND \$648 \$1064 \$1704 \$1587 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$4998 VPWR \$1735 VPWR VGND \$1384 \$1438 \$1679 VGND sky130_fd_sc_hd__or3_1
X$4999 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5000 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5001 VPWR \$1448 \$1736 \$1415 VPWR VGND \$1322 \$1705 VGND
+ sky130_fd_sc_hd__or4_1
X$5002 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5003 VGND \$1736 \$1811 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$5004 VPWR VGND VPWR \$1679 \$1705 VGND sky130_fd_sc_hd__inv_2
X$5005 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5008 VPWR \$1797 VPWR VGND \$1346 \$1662 VGND sky130_fd_sc_hd__or2_2
X$5009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5010 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5011 VPWR \$1631 VPWR VGND \$1766 VGND sky130_fd_sc_hd__buf_4
X$5012 VGND \$516 \$1707 \$1273 \$1708 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5013 VPWR VGND \$1680 \$542 \$1664 \$1641 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5014 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5015 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5016 VPWR \$1759 VGND VPWR \$1709 \$1363 \$1721 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$5017 VGND \$1709 \$411 \$1651 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5018 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5019 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5022 VGND \$516 \$1738 \$1273 \$1737 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5024 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5025 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5026 VGND \$1748 sram_ro_data[20] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$5027 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5028 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5030 VGND \$1762 \$1770 \$1376 \$1749 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$5031 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5032 VPWR \$1762 VGND VPWR \$1723 VGND sky130_fd_sc_hd__clkbuf_1
X$5033 VPWR \$1740 VGND VPWR \$1685 VGND sky130_fd_sc_hd__clkbuf_1
X$5034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5038 VPWR \$1742 VGND VPWR \$1689 VGND sky130_fd_sc_hd__clkbuf_1
X$5039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5041 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5044 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5045 VGND \$856 \$1772 \$1750 \$1751 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5047 VPWR VGND \$1815 VPWR \$1726 VGND sky130_fd_sc_hd__buf_2
X$5048 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5050 VGND \$463 \$1370 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5051 VPWR VGND \$1752 \$183 \$1728 \$1727 \$1774 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5055 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5057 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5058 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5059 VPWR \$1753 VGND VPWR \$1637 \$1776 \$815 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$5060 VGND \$1764 \$1753 \$1675 \$1715 \$1754 \$1007 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5062 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5063 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5065 VPWR \$1454 VGND VPWR \$1763 \$1034 VGND sky130_fd_sc_hd__or2_4
X$5066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5067 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5068 VGND \$1745 \$1693 \$1755 \$1125 \$1556 \$2013 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5069 VPWR VGND VPWR \$1640 \$1756 \$1765 \$1732 \$1745 VGND
+ sky130_fd_sc_hd__and4_1
X$5070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5071 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5072 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5076 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5077 VPWR VGND \$1572 \$183 \$1757 \$1794 \$1592 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5079 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5080 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5086 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5087 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5088 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5089 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5090 VPWR \$1704 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5092 VPWR \$1747 VPWR VGND \$1663 \$1746 \$1766 VGND sky130_fd_sc_hd__or3_1
X$5093 VGND \$1747 \$1743 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$5094 VGND \$1758 \$1776 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$5095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5096 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5097 VPWR \$1746 VPWR VGND \$1649 \$1532 VGND sky130_fd_sc_hd__or2_2
X$5098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5099 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5101 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5102 VPWR VGND VPWR \$1680 \$1681 VGND sky130_fd_sc_hd__inv_2
X$5103 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5104 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5105 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5107 VGND \$516 \$1721 \$1273 \$1759 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5108 VGND \$358 \$1273 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5109 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5110 VPWR \$1737 VGND VPWR \$1710 \$1363 \$1738 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$5111 VPWR VGND mgmt_gpio_oeb[4] VPWR \$1760 VGND sky130_fd_sc_hd__buf_2
X$5112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5114 VPWR \$1803 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5115 VPWR \$1767 VGND VPWR \$1803 VGND sky130_fd_sc_hd__clkbuf_1
X$5116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5117 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5119 VGND \$4776 \$4651 \$5104 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$5120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5121 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5122 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5123 VPWR \$5146 VGND VPWR \$4816 \$5076 \$907 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$5124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5126 VGND \$5154 \$1963 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$5127 VPWR \$5124 VGND VPWR \$4113 \$5089 VGND sky130_fd_sc_hd__or2b_2
X$5128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5129 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5130 VGND \$5110 \$3439 \$4576 VPWR VPWR VGND sky130_fd_sc_hd__nor2_4
X$5131 VPWR \$4476 VPWR VGND \$5110 \$5111 VGND sky130_fd_sc_hd__or2_2
X$5132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5133 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5134 VPWR \$4833 \$5091 \$4854 VPWR VGND \$5111 \$5090 VGND
+ sky130_fd_sc_hd__or4_1
X$5135 VPWR \$5093 VGND \$4476 \$5148 VPWR VGND sky130_fd_sc_hd__or2_1
X$5136 VPWR VGND \$4895 VPWR \$5112 VGND sky130_fd_sc_hd__clkbuf_4
X$5137 VPWR \$5105 VGND \$2552 \$4623 VPWR VGND sky130_fd_sc_hd__or2_1
X$5138 VPWR \$4777 VPWR VGND \$5113 \$4800 VGND sky130_fd_sc_hd__or2_2
X$5139 VPWR VGND \$4895 VPWR \$5106 \$2552 VGND sky130_fd_sc_hd__nor2_2
X$5140 VPWR \$5114 VPWR VGND \$5092 \$5105 VGND sky130_fd_sc_hd__nand2_1
X$5141 VPWR VPWR \$4623 VGND \$2996 \$5125 \$5114 VGND sky130_fd_sc_hd__o21bai_1
X$5142 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5143 VPWR \$5126 VGND \$4866 \$5125 VPWR VGND sky130_fd_sc_hd__or2_1
X$5144 VPWR VGND \$2996 VPWR \$4737 \$4953 VGND sky130_fd_sc_hd__nor2_2
X$5145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5146 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5149 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5151 VPWR VPWR \$5107 VGND \$5115 \$1369 \$4934 \$5033 VGND
+ sky130_fd_sc_hd__a211o_1
X$5152 VPWR \$5033 VGND \$1712 \$5116 VPWR VGND sky130_fd_sc_hd__or2_1
X$5153 VPWR \$4933 \$5116 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5154 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5157 VGND \$2777 \$5127 \$4811 \$5117 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5158 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5159 VPWR \$1557 \$5127 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$5160 VPWR VGND \$5118 \$3694 \$5064 \$5096 \$5080 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5162 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5163 VGND \$3694 \$542 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$5164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5166 VPWR VGND \$5081 VPWR \$5119 VGND sky130_fd_sc_hd__clkbuf_4
X$5167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5170 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5172 VGND \$4761 \$5066 \$4994 \$5128 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5173 VGND \$4761 \$5099 \$4994 \$5098 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5174 VPWR \$2854 \$5099 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$5175 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5176 VPWR VGND \$5044 \$4023 \$5083 \$5129 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5179 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5180 VPWR VGND \$4905 \$386 \$5085 \$5130 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5182 VPWR VGND \$5005 \$354 \$5108 \$5131 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5184 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5185 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5189 VPWR VGND \$4905 \$411 \$5120 \$5132 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5190 VPWR VGND \$5120 \$1423 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$5191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5192 VPWR VGND \$4905 \$354 \$5087 \$5133 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5193 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5194 VGND \$4764 \$5087 \$5006 \$5133 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5195 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5197 VGND \$4764 \$5102 \$4828 \$5101 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5198 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5199 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5200 VPWR VGND \$5046 \$411 \$5109 \$5135 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5201 VPWR VGND VPWR \$3825 \$5109 VGND sky130_fd_sc_hd__inv_2
X$5202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5203 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5204 VGND \$4764 \$5068 \$4828 \$5103 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5205 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5206 VPWR \$5137 VGND VPWR \$5121 \$4492 \$5122 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$5207 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5208 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5209 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5212 VGND \$5136 mgmt_gpio_out[15] \$2880 VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_2
X$5213 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5216 VPWR VGND wb_dat_o[25] VPWR \$5145 VGND sky130_fd_sc_hd__buf_2
X$5217 VPWR \$5153 VGND VPWR \$4862 \$5076 \$1829 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$5218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5219 VGND \$4816 \$4651 \$5146 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$5220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5221 VGND \$5138 \$1998 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$5222 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5223 VPWR \$5025 \$5138 \$4917 VPWR VGND \$4941 \$5147 VGND
+ sky130_fd_sc_hd__or4_1
X$5224 VPWR \$5111 VPWR VGND \$5089 \$5124 VGND sky130_fd_sc_hd__nand2_1
X$5225 VPWR \$4396 VPWR VGND \$4576 \$5139 VGND sky130_fd_sc_hd__or2_2
X$5226 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5227 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5228 VPWR \$4864 \$5112 \$4854 VPWR VGND \$5111 \$5148 VGND
+ sky130_fd_sc_hd__or4_1
X$5229 VPWR \$5140 VPWR VGND \$5111 \$5139 \$5148 VGND sky130_fd_sc_hd__or3_1
X$5230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5231 VPWR VGND \$4623 VPWR \$5140 VGND sky130_fd_sc_hd__buf_2
X$5232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5233 VPWR VGND VPWR \$5113 \$5105 VGND sky130_fd_sc_hd__inv_2
X$5234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5235 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5236 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5238 VPWR \$5141 VGND \$5126 VPWR \$5106 VGND sky130_fd_sc_hd__nor2_1
X$5239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5242 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5244 VGND \$3507 \$5149 VPWR \$1712 VPWR VGND sky130_fd_sc_hd__nand2_8
X$5245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5246 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5248 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5249 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5250 VPWR VGND \$5192 \$184 \$5127 \$5117 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5251 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5252 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5253 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5254 VPWR VGND \$5097 \$3711 \$5158 \$5157 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5255 VPWR \$3897 \$5156 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5257 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5258 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5259 VPWR VGND VPWR \$3417 \$5158 VGND sky130_fd_sc_hd__inv_2
X$5260 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5261 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5265 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5267 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5268 VGND \$4761 \$5083 \$4850 \$5129 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5269 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5270 VPWR VGND \$5044 \$4774 \$5150 \$5142 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5271 VPWR \$3886 \$5150 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5273 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5274 VGND \$4353 \$5085 \$4850 \$5130 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5275 VGND \$4764 \$5108 \$4850 \$5131 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5277 VPWR \$4058 \$5151 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5280 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5282 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5283 VGND \$4764 \$5120 \$5006 \$5132 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5285 VPWR VGND \$4905 \$542 \$5160 \$5143 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5286 VGND \$3952 \$5006 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5287 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5288 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5291 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5292 VGND \$4764 \$5109 \$4828 \$5135 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5293 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5294 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5295 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5296 VGND \$4764 \$5122 \$4828 \$5137 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5297 VGND \$5121 \$354 \$5161 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5300 VGND \$5144 \$1594 \$5162 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5302 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5306 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5307 VPWR \$1068 VPWR VGND \$1091 VGND sky130_fd_sc_hd__buf_4
X$5308 VPWR \$1111 VGND VPWR sram_ro_data[8] VGND sky130_fd_sc_hd__clkbuf_1
X$5309 VPWR \$1112 VGND VPWR sram_ro_data[9] VGND sky130_fd_sc_hd__clkbuf_1
X$5310 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5312 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5313 VPWR \$1102 VGND \$1092 VPWR \$918 VGND sky130_fd_sc_hd__or2b_1
X$5314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5318 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5319 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5322 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5323 VPWR \$1085 VPWR VGND \$1002 \$986 VGND sky130_fd_sc_hd__nand2_1
X$5324 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5325 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5326 VPWR VGND VPWR \$381 \$1086 VGND sky130_fd_sc_hd__inv_4
X$5327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5331 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5332 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5333 VGND \$856 \$1094 \$891 \$1095 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5335 VGND \$1113 \$1096 \$1103 \$1114 \$840 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$5336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5337 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5338 VGND \$463 \$922 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5341 VPWR VGND VPWR \$1115 \$1005 VGND sky130_fd_sc_hd__inv_2
X$5342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5343 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5344 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5347 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5348 VGND \$1104 \$1123 \$870 \$848 \$1103 \$1031 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5351 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5354 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5355 VPWR \$1105 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5356 VGND \$1117 \$753 \$365 \$1105 \$1116 \$1097 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$5357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5358 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5359 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5360 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5362 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5363 VPWR \$920 \$1035 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5365 VGND \$358 \$771 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5366 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5367 VPWR \$1118 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5368 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5369 VGND \$838 \$949 \$1107 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5371 VPWR \$1107 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5372 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5374 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5375 VGND \$1180 \$1106 \$620 \$379 \$433 \$217 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5380 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5383 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5387 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5392 VPWR VGND VPWR \$1110 \$1109 VGND sky130_fd_sc_hd__inv_2
X$5393 VGND \$1108 \$745 \$1120 \$1110 \$1012 VPWR VPWR VGND
+ sky130_fd_sc_hd__a22o_2
X$5394 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5395 VPWR VGND VPWR \$914 \$745 VGND sky130_fd_sc_hd__inv_2
X$5396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5397 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5400 VGND \$516 \$997 \$541 \$1013 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5405 VGND \$1131 sram_ro_data[10] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$5406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5407 VGND \$1143 \$945 \$1132 \$918 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5410 VPWR \$1144 VGND \$733 \$790 VPWR VGND sky130_fd_sc_hd__or2_1
X$5411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5412 VGND \$574 \$1122 \$1014 \$1069 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$5413 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5414 VGND \$1122 \$1015 \$790 \$1055 VPWR VPWR VGND sky130_fd_sc_hd__o21ai_4
X$5415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5419 VPWR VGND VPWR \$1145 \$1085 VGND sky130_fd_sc_hd__inv_2
X$5420 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5425 VPWR VGND \$1087 \$200 \$1146 \$1147 \$1088 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5426 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5427 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5428 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5429 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5433 VPWR \$1148 VGND VPWR \$1133 VGND sky130_fd_sc_hd__clkbuf_1
X$5434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5435 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5436 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5439 VPWR \$1149 VGND \$1116 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$5440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5441 VPWR \$1124 VGND VPWR \$338 \$320 \$1007 \$1116 VGND
+ sky130_fd_sc_hd__o22a_1
X$5442 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5444 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5445 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5446 VPWR \$1150 VGND VPWR \$1020 \$520 \$1232 \$1218 VGND
+ sky130_fd_sc_hd__o22a_1
X$5447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5449 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5450 VPWR \$1134 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5451 VPWR \$1106 VGND VPWR \$615 \$1103 \$1134 \$1125 VGND
+ sky130_fd_sc_hd__o22a_1
X$5452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5453 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5454 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5455 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5456 VGND \$1152 \$1151 \$605 \$1126 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5458 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5460 VPWR VGND \$990 \$200 \$1153 \$1154 \$991 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5461 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5462 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5465 VPWR VGND VPWR \$1155 \$949 VGND sky130_fd_sc_hd__inv_2
X$5466 VPWR \$1090 VGND VPWR \$1118 VGND sky130_fd_sc_hd__clkbuf_1
X$5467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5468 VPWR \$1127 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5469 VGND \$1119 \$949 \$1127 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5470 VGND \$1156 \$1135 \$259 \$326 \$1466 \$1099 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5472 VPWR \$1099 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5473 VPWR \$1157 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5474 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5475 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5477 VGND \$1136 \$578 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$5478 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5479 VGND \$516 \$1172 \$993 \$1158 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$5480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5481 VGND \$1159 \$1137 \$1128 \$1011 \$1138 VPWR VPWR VGND
+ sky130_fd_sc_hd__o31a_1
X$5482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5483 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5484 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5486 VGND \$516 \$1129 \$993 \$1160 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5488 VPWR \$1020 \$1139 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5490 VGND \$1161 \$914 \$1129 \$1140 \$1141 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$5491 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5492 VGND \$1108 \$1084 \$1109 \$1142 \$1184 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22ai_2
X$5493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5494 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5495 VGND \$516 \$745 \$466 \$1120 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$5496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5498 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5499 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5500 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5502 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5503 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5504 VPWR \$225 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5505 VPWR \$226 VGND \$235 VPWR \$236 VGND sky130_fd_sc_hd__or2b_1
X$5506 VPWR VGND sram_ro_addr[2] VPWR \$227 VGND sky130_fd_sc_hd__buf_2
X$5507 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5510 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5511 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5513 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5517 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5518 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5519 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5522 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5523 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5525 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5526 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5528 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5529 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5531 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5532 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5534 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5535 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5536 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5537 VGND \$206 \$223 \$243 \$232 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5539 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5541 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5542 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5543 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5544 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5545 VGND \$206 \$248 \$246 \$247 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5546 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5548 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5549 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5552 VGND \$206 \$222 \$246 \$250 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5553 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5554 VGND \$266 \$233 \$251 \$289 \$252 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$5555 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5556 VGND \$206 \$268 \$254 \$224 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5557 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5559 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5560 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5563 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5565 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5566 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5567 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5568 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5569 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5570 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5571 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5572 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5574 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5576 VPWR \$228 VGND VPWR \$302 VGND sky130_fd_sc_hd__clkbuf_1
X$5577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5578 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5580 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5581 VPWR \$238 VGND VPWR \$280 VGND sky130_fd_sc_hd__clkbuf_1
X$5582 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5584 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5585 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5587 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5588 VPWR VGND VPWR \$202 \$195 VGND sky130_fd_sc_hd__inv_2
X$5589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5590 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5591 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5592 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5594 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5595 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5598 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5602 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5604 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5605 VPWR \$229 \$230 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5608 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5610 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5611 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5613 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5615 VPWR \$287 VGND VPWR \$244 \$188 \$214 \$420 VGND sky130_fd_sc_hd__o22a_1
X$5616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5617 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5618 VPWR VGND \$271 \$294 \$223 \$232 \$288 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5620 VPWR VGND VPWR \$271 \$288 VGND sky130_fd_sc_hd__inv_2
X$5621 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5622 VPWR VGND \$271 \$200 \$296 \$209 \$288 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5624 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5625 VPWR \$1135 VGND VPWR \$245 \$188 \$256 \$456 VGND
+ sky130_fd_sc_hd__o22a_1
X$5626 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5627 VPWR \$278 VGND VPWR \$261 \$326 \$263 \$188 VGND sky130_fd_sc_hd__o22a_1
X$5628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5629 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5630 VPWR \$297 VGND VPWR \$210 \$433 \$191 \$755 VGND sky130_fd_sc_hd__o22a_1
X$5631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5632 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5633 VGND \$247 \$289 \$248 \$422 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$5634 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5635 VGND \$298 \$289 \$290 \$272 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$5636 VGND \$206 \$323 \$246 \$299 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5637 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5639 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5640 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5641 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5642 VGND \$206 \$252 \$246 \$266 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5644 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5645 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5646 VPWR VGND \$291 \$1179 \$300 \$279 \$292 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5647 VGND \$206 \$300 \$254 \$279 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$5648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5649 VPWR \$269 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5651 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5652 VPWR \$269 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5654 VPWR \$1171 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5655 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5657 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5658 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5659 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5660 VPWR VGND VPWR \$638 \$622 VGND sky130_fd_sc_hd__inv_2
X$5661 VPWR \$622 VGND VPWR sram_ro_data[0] VGND sky130_fd_sc_hd__clkbuf_1
X$5662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5663 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5665 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5666 VPWR \$629 VGND VPWR \$583 VGND sky130_fd_sc_hd__clkbuf_1
X$5667 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5668 VPWR \$596 VGND VPWR \$623 \$428 \$597 \$513 VGND sky130_fd_sc_hd__o22a_1
X$5669 VGND \$639 \$513 \$382 \$481 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$5670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5671 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5672 VPWR \$574 \$623 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5675 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5676 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5677 VPWR \$613 VGND VPWR \$586 VGND sky130_fd_sc_hd__clkbuf_1
X$5678 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5679 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5680 VGND \$655 \$555 \$237 \$614 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5681 VGND \$655 \$193 \$237 \$630 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$5682 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5683 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5684 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5688 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5689 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5693 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5694 VPWR VGND \$514 \$293 \$624 \$642 \$515 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5696 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5697 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5698 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5700 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5701 VGND \$516 \$603 \$196 \$625 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5702 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5703 VPWR \$631 \$603 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$5704 VGND \$516 \$604 \$196 \$632 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5706 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5708 VPWR VGND \$567 \$294 \$626 \$649 \$568 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5712 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5713 VPWR VGND \$627 \$281 \$617 \$606 \$607 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5714 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5715 VPWR VGND VPWR \$627 \$607 VGND sky130_fd_sc_hd__inv_2
X$5716 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5717 VGND \$516 \$608 \$243 \$618 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5719 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5720 VPWR VGND \$417 \$200 \$628 \$643 \$434 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5722 VGND \$644 \$223 \$662 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5723 VPWR VGND VPWR \$645 \$296 VGND sky130_fd_sc_hd__inv_2
X$5724 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5726 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5727 VGND \$633 \$296 \$619 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5728 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5729 VGND \$358 \$435 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$5730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5732 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5733 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5734 VGND \$532 \$593 \$671 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5735 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5736 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5737 VGND \$516 \$610 \$466 \$634 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5738 VGND \$634 \$289 \$610 \$647 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$5739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5740 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5741 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5743 VGND \$594 \$591 \$636 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5744 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5745 VPWR VGND VPWR \$289 \$612 VGND sky130_fd_sc_hd__inv_4
X$5746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5748 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5750 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5752 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5753 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5754 VPWR \$648 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5755 VPWR VGND mgmt_gpio_oeb[0] VPWR \$648 VGND sky130_fd_sc_hd__buf_2
X$5756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5758 VPWR \$653 VGND VPWR sram_ro_data[1] VGND sky130_fd_sc_hd__clkbuf_1
X$5759 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5763 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5764 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5770 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5771 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5772 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5773 VPWR VGND \$443 \$183 \$193 \$630 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5776 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5777 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5778 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5779 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5780 VGND \$655 \$641 \$241 \$656 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5781 VGND \$655 \$624 \$241 \$642 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5782 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5784 VPWR VGND \$514 \$200 \$658 \$657 \$515 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5786 VGND \$655 \$660 \$196 \$659 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5789 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5790 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5793 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5795 VGND \$516 \$626 \$605 \$649 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5796 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5799 VPWR VGND \$617 \$661 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$5800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5801 VPWR VGND \$608 \$646 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$5802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5804 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5806 VPWR \$662 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5808 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5809 VPWR \$662 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5811 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5812 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5813 VPWR VGND \$417 \$411 \$650 \$663 \$434 VPWR VGND sky130_fd_sc_hd__a22o_1
X$5814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5815 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5818 VGND \$516 \$593 \$466 \$651 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5819 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5820 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5821 VGND \$664 \$690 \$691 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5823 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5824 VGND \$647 \$665 \$664 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5825 VGND \$516 \$665 \$541 \$666 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5827 VPWR VGND VPWR \$289 \$611 VGND sky130_fd_sc_hd__inv_4
X$5828 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5829 VGND \$595 \$668 \$667 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$5830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5832 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5834 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5835 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5836 VGND \$206 \$571 \$246 \$652 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5837 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5838 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5841 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5843 VPWR VGND VPWR \$2485 \$1748 VGND sky130_fd_sc_hd__inv_2
X$5844 VPWR \$2423 VGND VPWR sram_ro_data[31] VGND sky130_fd_sc_hd__clkbuf_1
X$5845 VPWR \$2520 VGND VPWR \$2510 VGND sky130_fd_sc_hd__clkbuf_1
X$5846 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5847 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5848 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5851 VPWR \$2438 \$2437 VGND \$2487 VPWR \$2486 \$2512 VGND
+ sky130_fd_sc_hd__or4_2
X$5852 VPWR \$2513 \$2469 \$2521 VPWR VGND \$2468 \$2487 VGND
+ sky130_fd_sc_hd__or4_1
X$5853 VPWR \$2487 VGND \$2511 VPWR \$2514 VGND sky130_fd_sc_hd__nor2_1
X$5854 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5855 VPWR \$2353 VGND \$2472 VPWR \$2514 VGND sky130_fd_sc_hd__nor2_1
X$5856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5858 VPWR VGND VPWR \$2412 \$2453 VGND sky130_fd_sc_hd__inv_2
X$5859 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5860 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5861 VPWR VGND \$2472 \$2471 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$5862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5863 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5864 VPWR \$2393 VGND \$2511 VPWR \$2488 VGND sky130_fd_sc_hd__nor2_1
X$5865 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5866 VPWR \$2394 VGND \$2472 VPWR \$2488 VGND sky130_fd_sc_hd__nor2_1
X$5867 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5870 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5871 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5872 VPWR VGND \$1771 \$294 \$2490 \$2523 \$1815 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5874 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5875 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5876 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5879 VGND \$856 \$2455 \$1861 \$2491 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5880 VGND \$856 \$2473 \$1861 \$2492 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5881 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5882 VGND \$2280 \$2475 \$2522 \$2358 \$2274 \$2515 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5883 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5884 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5886 VGND \$2494 \$2493 \$1163 \$2525 \$2458 \$2516 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5887 VPWR \$2493 VGND VPWR \$1950 \$2456 \$2281 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$5888 VPWR VGND VPWR \$2526 \$2542 \$2494 \$2543 \$2370 VGND
+ sky130_fd_sc_hd__and4_1
X$5889 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5890 VPWR \$2527 VGND VPWR \$2457 \$1966 \$2176 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$5891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5892 VGND \$2496 \$1019 \$2005 \$2517 \$2300 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$5893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5894 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5895 VGND \$2526 \$2546 \$2496 \$2318 VPWR \$487 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$5896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5897 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5898 VGND \$2528 \$2271 \$2498 \$2162 \$859 \$1330 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5901 VGND \$2687 \$2852 \$2499 \$2501 VPWR \$662 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$5902 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5903 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5904 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5905 VGND \$2566 \$529 \$2502 \$1839 \$1507 \$796 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5908 VPWR \$2529 VGND VPWR \$861 \$2045 \$2503 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$5909 VPWR \$2480 VGND VPWR \$2498 \$1967 \$2518 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$5910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5911 VGND \$2530 \$2505 \$2460 \$2065 \$2046 \$2503 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5912 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5913 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5915 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5916 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5917 VPWR \$2506 VPWR VGND \$1438 \$1360 \$1679 VGND sky130_fd_sc_hd__or3_1
X$5918 VGND \$2506 \$2456 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$5919 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5920 VPWR \$1448 \$2532 \$1415 VPWR VGND \$1384 \$1679 VGND
+ sky130_fd_sc_hd__or4_1
X$5921 VPWR \$2507 VPWR VGND \$1322 \$1449 \$1705 VGND sky130_fd_sc_hd__or3_1
X$5922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5923 VPWR \$2533 VPWR VGND \$1322 \$1438 \$1679 VGND sky130_fd_sc_hd__or3_1
X$5924 VPWR \$1448 \$2534 \$1415 VPWR VGND \$1322 \$1679 VGND
+ sky130_fd_sc_hd__or4_1
X$5925 VGND \$2519 \$2559 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$5926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5928 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5929 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5930 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5933 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5934 VPWR VGND \$2127 \$184 \$2466 \$2484 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5935 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5938 VGND \$2535 \$2403 mgmt_gpio_out[6] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$5939 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5940 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5941 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5942 VPWR \$2550 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5943 VPWR \$2550 \$2510 VPWR \$1587 VGND VGND sky130_fd_sc_hd__and2_1
X$5944 VGND \$2233 \$2537 \$2119 \$2388 \$2570 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$5945 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5947 VPWR VGND VPWR \$2511 \$2390 VGND sky130_fd_sc_hd__inv_4
X$5948 VPWR \$2512 VPWR VGND \$2521 \$2436 \$2624 VGND sky130_fd_sc_hd__or3_1
X$5949 VPWR \$2468 VGND \$2514 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$5950 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5951 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5953 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5954 VPWR \$2391 VGND \$2453 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$5955 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5959 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5961 VPWR \$2538 VGND \$2553 \$2489 VPWR VGND sky130_fd_sc_hd__or2_1
X$5962 VGND \$856 \$2555 \$1750 \$2554 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$5963 VGND \$856 \$2490 \$2556 \$2523 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$5964 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5965 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5966 VPWR VGND \$2321 \$281 \$2557 \$2572 \$2322 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5967 VPWR VGND \$2321 \$294 \$2558 \$2573 \$2322 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$5968 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5969 VPWR \$2574 VGND VPWR \$1722 \$1554 \$2382 \$923 VGND
+ sky130_fd_sc_hd__o22a_1
X$5970 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5971 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5973 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5974 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5975 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5976 VPWR VGND VPWR \$2457 \$2473 VGND sky130_fd_sc_hd__inv_2
X$5977 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$5978 VPWR \$2575 VGND VPWR \$1256 \$2135 \$2292 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$5979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5981 VPWR \$2577 VGND VPWR \$1081 \$2559 \$2539 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$5982 VGND \$2543 \$2577 \$2342 \$2750 \$2541 \$756 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5983 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5984 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$5987 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5988 VGND \$2546 \$2560 \$2515 \$2544 \$2545 \$2298 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$5990 VPWR \$1676 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$5991 VGND \$2563 \$2345 \$2457 \$2190 \$1676 \$2561 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5992 VGND \$2580 \$2562 \$2292 \$1729 \$2497 \$2518 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$5993 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$5994 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$5995 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$5996 VPWR \$1420 VGND VPWR \$2447 \$1571 VGND sky130_fd_sc_hd__or2_4
X$5997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$5998 VPWR VGND VPWR \$2585 \$2564 \$2578 \$2584 \$2583 VGND
+ sky130_fd_sc_hd__and4_1
X$5999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6000 VPWR VGND VPWR \$2564 \$2566 \$2586 \$2565 \$2429 VGND
+ sky130_fd_sc_hd__and4_1
X$6001 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6002 VPWR \$2547 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$6003 VGND \$2586 \$2303 \$2460 \$1867 \$2614 \$2547 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6004 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6005 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6006 VGND \$2588 \$2399 \$2460 \$2047 \$2048 \$2587 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6008 VGND \$2567 \$2568 \$2589 \$2530 VPWR \$968 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$6009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6010 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6011 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6013 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6014 VGND \$2569 \$2750 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6016 VGND \$2508 \$2541 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6017 VPWR \$1448 \$2591 \$1415 VPWR VGND \$1882 \$1679 VGND
+ sky130_fd_sc_hd__or4_1
X$6018 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6019 VGND \$2533 \$2540 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6023 VGND \$2462 \$2544 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$6024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6025 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6027 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6029 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6031 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6032 VGND \$2535 \$2620 \$1721 \$2551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6033 VPWR \$2548 \$2466 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6036 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6037 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6038 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6043 VPWR \$1350 \$1366 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6044 VPWR \$1366 VGND VPWR sram_ro_data[13] VGND sky130_fd_sc_hd__clkbuf_1
X$6045 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6046 VPWR \$1247 \$1367 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6051 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6052 VPWR \$1375 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$6053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6057 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6058 VPWR \$1377 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$6059 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6060 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6062 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6063 VGND \$1336 \$1162 \$1368 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6064 VGND \$1352 \$1337 \$1376 \$1314 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6066 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6067 VGND \$1369 \$1230 \$2070 \$1353 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$6068 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6069 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6070 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6071 VGND \$1378 \$1460 \$1354 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6072 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6073 VGND \$856 \$1388 \$1370 \$1355 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6076 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6077 VPWR VGND VPWR \$1299 \$856 VGND sky130_fd_sc_hd__inv_2
X$6078 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6079 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6080 VGND \$1299 \$1341 \$565 VPWR VPWR VGND sky130_fd_sc_hd__nor2_8
X$6081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6082 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6083 VPWR \$1356 VGND VPWR \$816 \$1342 VGND sky130_fd_sc_hd__or2_4
X$6084 VPWR \$1356 VGND VPWR \$1103 \$1248 VGND sky130_fd_sc_hd__or2_4
X$6085 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6086 VGND \$1318 \$1401 \$1379 \$1389 \$1317 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6087 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6088 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6090 VGND \$1353 \$1283 \$1317 \$1412 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6092 VGND \$1372 \$1371 \$1192 \$1271 \$816 \$1115 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6093 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6094 VPWR \$1258 VGND VPWR \$1198 \$1342 VGND sky130_fd_sc_hd__or2_4
X$6095 VPWR VGND VPWR \$1381 \$1316 \$1372 \$1104 \$1380 VGND
+ sky130_fd_sc_hd__and4_1
X$6096 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6097 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6099 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6100 VGND \$655 \$1357 \$605 \$1319 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6101 VGND \$1382 \$1331 \$1373 \$1089 \$686 \$936 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6102 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6103 VPWR VGND \$1178 \$183 \$1332 \$1343 \$1166 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6105 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6107 VPWR VGND \$990 \$281 \$1358 \$1403 \$991 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6108 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6110 VPWR VGND VPWR \$1383 \$1344 VGND sky130_fd_sc_hd__inv_2
X$6111 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6112 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6113 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6114 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6116 VPWR VGND \$1295 VPWR \$1359 VGND sky130_fd_sc_hd__buf_2
X$6117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6118 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6121 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6122 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6123 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6124 VPWR \$1137 VGND VPWR \$1384 \$1345 VGND sky130_fd_sc_hd__or2_4
X$6125 VPWR VGND VPWR \$1345 \$1138 VGND sky130_fd_sc_hd__inv_2
X$6126 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6127 VPWR VGND VPWR \$1361 \$1449 VGND sky130_fd_sc_hd__inv_2
X$6128 VGND \$1362 \$1011 \$1212 \$1361 \$1323 \$1374 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$6129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6130 VPWR VGND VPWR \$1346 \$1308 VGND sky130_fd_sc_hd__inv_2
X$6131 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6133 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6135 VGND \$516 \$1415 \$541 \$1392 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$6136 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6137 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6138 VPWR \$1407 VGND VPWR \$1364 \$1363 \$1354 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$6139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6140 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6141 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6143 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6144 VPWR VGND VPWR \$1365 \$1363 VGND sky130_fd_sc_hd__inv_2
X$6145 VGND \$358 \$1274 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$6146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6150 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6151 VPWR \$1395 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$6152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6154 VPWR \$1395 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$6155 VGND \$1409 \$1186 \$564 \$1396 \$780 \$1144 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$6156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6157 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6158 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6159 VGND \$1410 \$1385 \$1396 \$1014 \$574 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$6160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6162 VGND \$1416 \$1433 \$1376 \$1397 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$6163 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6164 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6165 VGND \$1145 \$1386 \$1162 \$1337 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$6166 VPWR \$1368 VGND \$1351 VPWR \$1386 VGND sky130_fd_sc_hd__nor2_1
X$6167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6168 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6170 VGND \$1387 \$1162 \$1337 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6171 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6172 VGND \$1369 \$1229 \$1398 \$1412 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$6173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6174 VGND \$1215 \$1385 \$1083 \$1315 VPWR VPWR VGND sky130_fd_sc_hd__o21ai_4
X$6175 VPWR VGND \$1399 \$293 \$1388 \$1355 \$1417 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6177 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6178 VGND \$856 \$1418 \$1370 \$1400 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6181 VGND \$484 \$1411 \$1248 \$1401 VPWR VPWR VGND sky130_fd_sc_hd__or3b_4
X$6182 VPWR \$1401 VGND VPWR \$686 \$1248 VGND sky130_fd_sc_hd__or2_4
X$6183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6184 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6185 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6186 VGND \$1389 \$1356 \$1317 \$1412 \$1379 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6187 VPWR \$1389 \$1353 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6188 VPWR \$1326 \$1379 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6189 VGND \$1412 \$1059 \$1326 \$1389 \$1328 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6190 VPWR \$1328 \$1317 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6192 VGND \$1353 \$1420 \$1317 \$1412 \$1379 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6193 VGND \$1318 \$1264 \$1379 \$1353 \$1317 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$6194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6195 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6198 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6199 VPWR \$1402 VGND VPWR \$1247 \$1297 \$403 \$420 VGND
+ sky130_fd_sc_hd__o22a_1
X$6200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6201 VPWR VPWR VGND \$966 \$1201 VGND sky130_fd_sc_hd__clkbuf_2
X$6202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6204 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6207 VPWR VGND VPWR \$1390 \$1357 VGND sky130_fd_sc_hd__inv_2
X$6208 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6209 VPWR VGND VPWR \$1080 \$1332 VGND sky130_fd_sc_hd__inv_2
X$6210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6212 VGND \$1152 \$1358 \$771 \$1403 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6213 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6214 VPWR VPWR VGND \$1404 \$991 VGND sky130_fd_sc_hd__clkbuf_2
X$6215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6217 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6220 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6222 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6223 VPWR VGND \$1170 \$294 \$1413 \$1391 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6225 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6226 VGND \$1128 \$1322 \$531 \$1705 VPWR VPWR VGND sky130_fd_sc_hd__nor3_4
X$6227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6228 VPWR \$1405 VGND \$1415 \$1374 VPWR VGND sky130_fd_sc_hd__or2_1
X$6229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6230 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6231 VPWR \$1405 VPWR VGND \$1128 VGND sky130_fd_sc_hd__buf_4
X$6232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6233 VPWR \$1562 VPWR VGND \$503 \$1406 \$1299 VGND sky130_fd_sc_hd__or3_2
X$6234 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6236 VPWR VGND \$672 \$1415 \$1414 \$1392 \$895 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6237 VPWR VGND VPWR \$1414 \$1415 VGND sky130_fd_sc_hd__inv_2
X$6238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6240 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6241 VGND \$516 \$1354 \$1273 \$1407 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$6242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6244 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6245 VGND \$1393 \$386 \$1275 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6247 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6250 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6252 VPWR \$2166 \$2153 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6253 VPWR VGND VPWR \$2091 \$2129 VGND sky130_fd_sc_hd__inv_2
X$6254 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6255 VPWR \$2167 VGND VPWR \$2210 VGND sky130_fd_sc_hd__clkbuf_1
X$6256 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6257 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6258 VPWR \$2168 VGND \$2154 \$1963 VPWR VGND sky130_fd_sc_hd__or2_1
X$6259 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6260 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6261 VGND \$2212 \$1960 \$2169 \$2155 \$2130 \$1897 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_4
X$6262 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6263 VPWR \$2132 VPWR VGND \$2188 \$2131 \$2025 VGND sky130_fd_sc_hd__or3_1
X$6264 VPWR \$1977 VPWR VGND \$1919 \$1933 \$2131 VGND sky130_fd_sc_hd__or3_1
X$6265 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6267 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6268 VGND \$2156 \$2171 \$2133 \$2170 \$2132 \$2172 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2111o_2
X$6269 VPWR VGND VPWR \$2172 \$2119 VGND sky130_fd_sc_hd__inv_2
X$6270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6271 VPWR \$2173 VGND \$2026 VPWR \$1962 VGND sky130_fd_sc_hd__nor2_1
X$6272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6275 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6276 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6279 VGND \$856 \$2134 \$1370 \$2157 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6280 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6281 VPWR \$2174 VGND VPWR \$506 \$456 \$2091 \$1556 VGND
+ sky130_fd_sc_hd__o22a_1
X$6282 VPWR VGND \$1752 \$293 \$2158 \$2175 \$1774 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6284 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6285 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6287 VPWR \$2176 \$2084 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6288 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6289 VPWR VGND VPWR \$2120 \$2106 VGND sky130_fd_sc_hd__inv_2
X$6290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6292 VPWR VGND VPWR \$1965 \$2071 VGND sky130_fd_sc_hd__inv_2
X$6293 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6294 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6295 VPWR \$2177 VGND VPWR \$1282 \$2135 \$2018 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$6296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6297 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6298 VGND \$2125 \$2159 \$601 \$785 \$2220 \$1325 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6299 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6300 VPWR VGND VPWR \$2137 \$2074 \$2105 \$2136 \$2178 VGND
+ sky130_fd_sc_hd__and4_1
X$6301 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6302 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6303 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6304 VGND \$2179 \$726 \$2005 \$2160 \$2140 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$6305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6306 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6307 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6309 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6310 VPWR \$2087 VGND VPWR \$784 \$2045 \$1080 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$6311 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6312 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6313 VGND \$2181 \$2174 \$1965 \$2190 \$2180 \$1915 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6315 VGND \$2182 \$1843 \$2161 \$2065 \$2046 \$1080 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6317 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6318 VGND \$2178 \$2112 \$2161 \$2047 \$2048 \$819 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6321 VGND \$2142 \$2141 \$758 \$379 \$2162 \$2163 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6322 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6323 VGND \$1152 \$2143 \$1627 \$2144 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6324 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6325 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6328 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6330 VPWR \$2183 VGND \$2080 \$1780 VPWR VGND sky130_fd_sc_hd__or2_1
X$6331 VPWR \$2164 VGND \$1813 \$1780 VPWR VGND sky130_fd_sc_hd__or2_1
X$6332 VPWR \$2184 VPWR VGND \$1814 \$1797 \$1766 VGND sky130_fd_sc_hd__or3_1
X$6333 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6334 VGND \$2147 \$785 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6335 VGND \$2148 \$2116 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6336 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6337 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6338 VGND \$2149 \$804 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$6339 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6340 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6341 VPWR VGND VPWR \$3005 \$2101 VGND sky130_fd_sc_hd__inv_2
X$6342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6344 VPWR VGND \$1680 \$184 \$2165 \$2150 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6346 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6347 VPWR VGND VPWR \$1823 \$2151 VGND sky130_fd_sc_hd__inv_2
X$6348 VGND \$1152 \$2151 \$2232 \$2185 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6349 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6352 VGND \$2068 \$2033 mgmt_gpio_out[5] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$6353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6355 VGND \$2167 \$2040 \$1376 \$2039 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$6356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6357 VGND \$2014 \$2168 \$2195 \$2211 \$2001 \$2194 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$6358 VGND \$2212 \$2195 \$2194 \$2119 \$2154 \$1962 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6359 VPWR VPWR \$2155 \$2188 \$2193 \$2187 \$2194 \$2119 VGND VGND
+ sky130_fd_sc_hd__o2111ai_1
X$6360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6361 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6364 VPWR \$2170 VGND \$2119 VPWR \$2002 VGND sky130_fd_sc_hd__nor2_1
X$6365 VPWR \$2196 VPWR VGND \$2041 \$1921 \$2170 VGND sky130_fd_sc_hd__or3_1
X$6366 VPWR \$2196 \$2189 VGND \$2133 VPWR \$2197 \$1978 VGND
+ sky130_fd_sc_hd__or4_2
X$6367 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6368 VPWR VPWR \$2223 VGND \$2172 \$2171 \$2104 \$2173 VGND
+ sky130_fd_sc_hd__a211o_1
X$6369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6370 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6371 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6372 VPWR \$2217 VGND \$2198 \$2059 VPWR VGND sky130_fd_sc_hd__or2_1
X$6373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6376 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6377 VPWR VGND \$1923 \$294 \$2199 \$2245 \$1924 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6380 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6382 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6383 VGND \$856 \$2158 \$1861 \$2175 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6387 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6389 VPWR \$1356 VGND VPWR \$2190 \$1571 VGND sky130_fd_sc_hd__or2_4
X$6390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6391 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6394 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6395 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6399 VGND \$2459 \$2200 \$2179 \$2182 VPWR \$512 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$6400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6403 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6405 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6406 VGND \$4238 \$2076 \$2190 \$2113 \$2161 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$6407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6409 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6411 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6413 VPWR VGND VPWR \$2161 \$2143 VGND sky130_fd_sc_hd__inv_2
X$6414 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6418 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6419 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6420 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6421 VPWR \$2201 VGND \$2080 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$6422 VGND \$2164 \$2358 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6424 VGND \$2184 \$2220 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6427 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6428 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6429 VPWR \$2202 VGND \$1531 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$6430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6431 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6432 VPWR \$1867 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$6433 VPWR \$2192 VGND \$1867 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$6434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6436 VPWR VGND \$1680 \$1171 \$2203 \$2204 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6437 VGND \$358 \$2937 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$6438 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6439 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6440 VPWR VGND \$2128 VPWR \$2192 VGND sky130_fd_sc_hd__buf_2
X$6441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6444 VPWR VGND \$2127 \$1179 \$2205 \$2206 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6445 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6446 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6447 VPWR VGND \$2127 \$542 \$2207 \$2208 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6450 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6454 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6455 VPWR VGND wb_dat_o[31] VPWR \$5403 VGND sky130_fd_sc_hd__buf_2
X$6456 VGND \$5024 \$5002 \$5374 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$6457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6458 VGND \$5001 \$5002 \$5395 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$6459 VPWR \$5395 VGND VPWR \$5001 \$5076 \$1975 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$6460 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6461 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6463 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6465 VGND \$4632 \$5404 \$2472 \$4474 \$5268 \$5326 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$6466 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6467 VPWR VGND \$5025 \$4930 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$6468 VPWR \$5268 VGND \$5405 \$2571 VPWR VGND sky130_fd_sc_hd__or2_1
X$6469 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6470 VPWR \$5281 \$4941 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$6471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6472 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6473 VGND \$5386 \$2741 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$6474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6475 VPWR \$5406 VPWR VGND \$5281 \$4930 \$4917 VGND sky130_fd_sc_hd__or3_1
X$6476 VPWR \$5405 VPWR \$5219 VGND VGND sky130_fd_sc_hd__clkinvlp_2
X$6477 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6478 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6479 VPWR \$5422 VGND VPWR \$4752 \$4892 VGND sky130_fd_sc_hd__or2b_2
X$6480 VPWR \$5359 VGND \$5147 \$5281 VPWR VGND sky130_fd_sc_hd__or2_1
X$6481 VPWR \$5396 VPWR VGND \$5025 \$4942 \$5359 VGND sky130_fd_sc_hd__or3_1
X$6482 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6483 VGND \$5396 \$2472 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$6484 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6485 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6486 VGND \$5375 \$2511 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6488 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6491 VPWR \$5336 VPWR VGND \$5303 \$5440 \$5348 VGND sky130_fd_sc_hd__or3_2
X$6492 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6495 VPWR \$5284 VGND \$2511 VPWR \$5415 VGND sky130_fd_sc_hd__nor2_1
X$6496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6500 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6503 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6506 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6507 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6511 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6513 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6518 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6519 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6520 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6521 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6522 VGND \$2777 \$5387 \$5165 \$5397 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6523 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6524 VPWR VGND \$5192 \$4023 \$5387 \$5397 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6526 VPWR \$1235 \$5387 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$6527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6528 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6529 VGND \$4761 \$5341 \$5165 \$5379 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6532 VGND \$4761 \$5380 \$5165 \$5381 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6534 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6535 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6536 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6538 VGND \$4761 \$5389 \$5408 \$5398 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$6539 VPWR VGND \$5388 \$184 \$5389 \$5398 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6540 VPWR VGND \$5390 VPWR \$5238 VGND sky130_fd_sc_hd__clkbuf_4
X$6541 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6542 VGND \$4761 \$5364 \$4994 \$5382 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6543 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6544 VPWR \$1134 \$5389 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$6545 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6547 VGND \$4374 \$4994 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$6548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6549 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6550 VGND \$4761 \$5365 \$4994 \$5409 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6552 VPWR VGND VPWR \$5252 \$5262 VGND sky130_fd_sc_hd__inv_2
X$6553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6554 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6555 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6558 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6559 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6561 VPWR VGND \$5332 \$1171 \$5331 \$5366 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6562 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6563 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6565 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6566 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6567 VGND \$4761 \$5368 \$5367 \$5402 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6568 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6569 VPWR VGND \$5332 \$386 \$5368 \$5402 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6573 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6575 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6576 VGND \$4761 \$5392 \$5369 \$5410 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6577 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6578 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6579 VPWR VGND VPWR \$3254 \$5392 VGND sky130_fd_sc_hd__inv_2
X$6580 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6582 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6583 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6586 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6587 VPWR VGND \$5332 \$354 \$5333 \$5383 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6588 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6591 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6592 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6593 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6594 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6595 VGND \$4764 \$5371 \$5334 \$5399 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6596 VPWR VGND \$5344 \$4774 \$5371 \$5399 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6599 VPWR VGND \$5344 \$184 \$5372 \$5384 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6600 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6601 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6603 VGND \$4764 \$5372 \$5334 \$5384 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6604 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6606 VGND \$4764 \$5385 \$5334 \$5400 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6607 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6608 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6609 VPWR VGND \$5345 \$3694 \$5385 \$5400 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6614 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6616 VPWR \$5411 VGND VPWR \$5401 \$4724 \$5413 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$6617 VGND \$5401 \$354 \$5299 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6618 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6619 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6621 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6622 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6628 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6629 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6630 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6631 VPWR VGND VPWR \$4609 \$5393 VGND sky130_fd_sc_hd__inv_2
X$6632 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6637 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6638 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6639 VPWR VGND VPWR \$778 \$767 VGND sky130_fd_sc_hd__inv_2
X$6640 VPWR VGND VPWR \$718 \$747 VGND sky130_fd_sc_hd__inv_4
X$6641 VPWR \$767 VGND VPWR sram_ro_data[3] VGND sky130_fd_sc_hd__clkbuf_1
X$6642 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6643 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6644 VPWR \$719 VGND VPWR \$738 VGND sky130_fd_sc_hd__clkbuf_1
X$6645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6646 VGND \$738 \$720 \$779 \$918 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6647 VGND \$779 \$780 \$768 \$564 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6649 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6651 VPWR VGND \$720 \$768 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$6652 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6653 VPWR \$597 VPWR VGND \$733 \$481 \$382 VGND sky130_fd_sc_hd__or3_2
X$6654 VGND \$781 \$597 \$382 \$481 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$6655 VPWR \$748 VGND \$439 VPWR \$481 VGND sky130_fd_sc_hd__nor2_1
X$6656 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6657 VPWR \$382 VPWR \$1079 VGND \$597 \$481 VGND sky130_fd_sc_hd__o21a_1
X$6658 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6659 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6660 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6661 VPWR \$750 VPWR VGND \$739 \$749 \$439 VGND sky130_fd_sc_hd__or3_1
X$6662 VPWR VGND VPWR \$739 \$597 VGND sky130_fd_sc_hd__inv_2
X$6663 VPWR VGND \$623 VPWR \$750 VGND sky130_fd_sc_hd__clkbuf_4
X$6664 VPWR VGND VPWR \$749 \$481 VGND sky130_fd_sc_hd__inv_2
X$6665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6666 VPWR \$739 \$740 \$790 VPWR VGND \$439 \$749 VGND sky130_fd_sc_hd__or4_1
X$6667 VGND \$751 \$673 \$721 \$1015 \$681 \$623 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$6668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6669 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6670 VPWR VGND VPWR \$721 \$682 VGND sky130_fd_sc_hd__inv_2
X$6671 VPWR VGND VPWR \$681 \$740 VGND sky130_fd_sc_hd__inv_2
X$6672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6673 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6674 VPWR VGND \$740 \$741 \$682 \$734 \$681 VPWR VGND sky130_fd_sc_hd__a22o_1
X$6675 VGND \$722 \$741 \$381 \$734 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$6676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6678 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6681 VGND \$655 \$227 \$237 \$752 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$6682 VPWR VGND \$443 \$200 \$227 \$752 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$6683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6685 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6688 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6689 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6691 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6693 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6694 VGND \$655 \$724 \$241 \$723 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6697 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6698 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6699 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6701 VPWR VGND VPWR \$769 \$724 VGND sky130_fd_sc_hd__inv_2
X$6702 VGND \$655 \$783 \$241 \$761 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6706 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6710 VPWR VPWR VGND \$742 \$515 VGND sky130_fd_sc_hd__clkbuf_2
X$6711 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6713 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6714 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6718 VPWR VGND \$602 \$294 \$743 \$735 \$674 VPWR VGND sky130_fd_sc_hd__a22o_1
X$6719 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6720 VGND \$655 \$743 \$196 \$735 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6722 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6724 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6725 VPWR VGND \$743 \$762 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$6726 VPWR \$727 VGND \$744 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$6727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6729 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6730 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6731 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6732 VGND \$655 \$728 \$605 \$736 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6733 VGND \$881 \$763 \$755 \$744 \$703 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$6734 VPWR \$784 \$528 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6735 VPWR \$770 \$728 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6736 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6737 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6738 VGND \$753 \$590 \$500 \$379 \$744 \$616 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$6739 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6740 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6742 VGND \$754 \$687 \$744 \$755 \$635 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$6743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6744 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6745 VPWR VGND VPWR \$756 \$729 VGND sky130_fd_sc_hd__inv_2
X$6746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6748 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6749 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6750 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6751 VGND \$516 \$737 \$771 \$757 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6752 VPWR VGND \$627 \$294 \$737 \$757 \$607 VPWR VGND sky130_fd_sc_hd__a22o_1
X$6753 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6754 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6755 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6756 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6757 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6758 VPWR VGND \$417 \$294 \$772 \$786 \$434 VPWR VGND sky130_fd_sc_hd__a22o_1
X$6759 VPWR VGND VPWR \$758 \$628 VGND sky130_fd_sc_hd__inv_2
X$6760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6762 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6763 VPWR VGND \$434 VPWR \$773 VGND sky130_fd_sc_hd__clkbuf_4
X$6764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6766 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6767 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6770 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6771 VPWR VGND VPWR \$713 \$714 VGND sky130_fd_sc_hd__inv_2
X$6772 VGND \$3655 \$764 \$755 \$774 \$848 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_4
X$6773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6775 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6778 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6779 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6781 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6783 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6784 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6785 VGND \$788 \$289 \$775 \$765 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$6786 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6788 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6789 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6793 VGND \$516 \$789 \$466 \$766 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6794 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6795 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6796 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6798 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6799 VPWR VGND VPWR \$289 \$715 VGND sky130_fd_sc_hd__inv_4
X$6800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6804 VPWR VGND VPWR \$289 \$716 VGND sky130_fd_sc_hd__inv_4
X$6805 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6806 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6808 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6809 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6810 VPWR VGND VPWR \$696 \$677 VGND sky130_fd_sc_hd__inv_2
X$6811 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6812 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6815 VPWR VGND VPWR \$717 \$984 VGND sky130_fd_sc_hd__inv_2
X$6816 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6817 VGND \$889 \$698 \$776 \$808 \$777 \$697 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$6818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6819 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6820 VGND \$206 \$759 \$246 \$746 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6821 VPWR VGND VPWR \$777 \$698 VGND sky130_fd_sc_hd__inv_2
X$6822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6823 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6828 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6829 VPWR VGND wb_dat_o[21] VPWR \$5001 VGND sky130_fd_sc_hd__buf_2
X$6830 VGND \$4950 \$4651 \$4976 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$6831 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6832 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6833 VGND \$4622 \$5002 \$5012 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$6834 VPWR \$4508 \$4509 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6835 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6836 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6837 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6840 VGND \$5013 \$1962 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$6841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6842 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6843 VPWR \$4951 VGND \$4394 \$4917 VPWR VGND sky130_fd_sc_hd__or2_1
X$6844 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6845 VGND \$5003 \$2742 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6846 VGND \$4977 \$2700 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$6847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6849 VPWR \$5025 \$4910 \$4986 VPWR VGND \$4698 \$4444 VGND
+ sky130_fd_sc_hd__or4_1
X$6850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6851 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6852 VPWR \$4987 VPWR VGND \$4864 \$4892 \$4757 VGND sky130_fd_sc_hd__or3_1
X$6853 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6856 VPWR \$4882 VGND \$4987 VPWR \$4394 VGND sky130_fd_sc_hd__nor2_1
X$6857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6858 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6859 VPWR \$5014 VGND \$5004 VPWR \$4855 VGND sky130_fd_sc_hd__nor2_1
X$6860 VGND \$4006 \$4326 \$4673 VPWR VPWR VGND sky130_fd_sc_hd__nor2_4
X$6861 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6862 VPWR VGND VPWR \$4912 \$4987 VGND sky130_fd_sc_hd__inv_2
X$6863 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6864 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6865 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6866 VPWR VPWR \$2742 VGND \$4623 \$4988 \$5015 VGND sky130_fd_sc_hd__o21bai_1
X$6867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6868 VPWR \$5016 VPWR VGND \$4267 \$4989 \$4988 VGND sky130_fd_sc_hd__or3_1
X$6869 VPWR VGND \$4882 VPWR \$4942 \$4978 \$4962 VGND sky130_fd_sc_hd__a21o_1
X$6870 VPWR \$4978 VGND \$5016 \$4326 VPWR VGND sky130_fd_sc_hd__or2_1
X$6871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6872 VPWR \$4989 VGND \$4895 VPWR \$2742 VGND sky130_fd_sc_hd__nor2_1
X$6873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6874 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6875 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6876 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6877 VPWR VPWR \$4953 VGND \$2700 \$4932 \$5060 VGND sky130_fd_sc_hd__o21ai_1
X$6878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6879 VPWR \$4964 VGND \$2700 VPWR \$4953 VGND sky130_fd_sc_hd__nor2_1
X$6880 VPWR \$5017 VGND \$4617 \$4990 VPWR VGND sky130_fd_sc_hd__or2_1
X$6881 VPWR \$4990 VGND \$4963 VPWR \$4964 VGND sky130_fd_sc_hd__nor2_1
X$6882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6883 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6884 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6886 VPWR \$5034 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$6887 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6888 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6889 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6890 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6892 VGND \$2777 \$4979 \$4811 \$4991 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6894 VPWR VGND \$4701 \$3694 \$4979 \$4991 \$4677 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6895 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6896 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6897 VPWR VGND \$4979 \$3129 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$6898 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6901 VPWR VGND \$4760 \$293 \$4955 \$4992 \$4717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6904 VGND \$4761 \$4944 \$4406 \$4965 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6906 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6907 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6908 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6909 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6910 VGND \$4761 \$4967 \$4813 \$4966 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6911 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6912 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6913 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6915 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6916 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6917 VGND \$4374 \$4813 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$6918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6919 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6920 VPWR VGND \$4654 \$354 \$4937 \$4968 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6921 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6924 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6925 VGND \$4761 \$4980 \$4813 \$4993 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6927 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6928 VPWR \$3937 \$4980 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6930 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6931 VPWR VGND \$5005 \$4023 \$4980 \$4993 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6932 VGND \$4353 \$4958 \$4994 \$4969 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6933 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6934 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6935 VGND \$4353 \$4981 \$4850 \$4995 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6937 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6938 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6939 VPWR \$4028 \$4981 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6940 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6941 VPWR VGND \$5005 \$1594 \$5020 \$5019 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6943 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6944 VPWR VGND VPWR \$2615 \$5020 VGND sky130_fd_sc_hd__inv_2
X$6945 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6946 VGND \$4353 \$4959 \$4850 \$4970 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$6947 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6949 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6950 VGND \$4764 \$4982 \$4850 \$4996 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6951 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6952 VPWR VGND \$5005 \$411 \$4982 \$4996 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6954 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6955 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6958 VPWR VGND \$4899 \$411 \$4938 \$4971 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$6960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6961 VGND \$4764 \$4960 \$4765 \$4972 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6963 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6966 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$6967 VPWR VGND \$4899 \$354 \$4983 \$4997 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6968 VGND \$4764 \$4983 \$5006 \$4997 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6969 VPWR VGND \$4900 VPWR \$4973 VGND sky130_fd_sc_hd__clkbuf_4
X$6970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6971 VPWR VGND VPWR \$4482 \$4983 VGND sky130_fd_sc_hd__inv_2
X$6972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6973 VPWR VGND VPWR \$4905 \$5100 VGND sky130_fd_sc_hd__inv_2
X$6974 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6975 VPWR VGND \$5035 VPWR \$4794 VGND sky130_fd_sc_hd__clkbuf_4
X$6976 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6977 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6978 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6979 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6980 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6981 VGND \$5007 \$4482 \$2614 \$4239 \$5008 \$3659 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$6982 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$6983 VPWR \$4017 \$5009 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$6984 VPWR VGND \$4998 VPWR \$4767 VGND sky130_fd_sc_hd__clkbuf_4
X$6985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6987 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6988 VPWR VGND VPWR \$4039 \$4984 VGND sky130_fd_sc_hd__inv_2
X$6989 VPWR VGND \$5046 \$386 \$4984 \$4999 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$6990 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$6991 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$6992 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6993 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6994 VPWR VGND VPWR \$5010 \$2900 VGND sky130_fd_sc_hd__inv_4
X$6995 VGND \$4764 \$5010 \$4828 \$5022 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$6996 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$6997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$6998 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$6999 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7000 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7002 VGND \$2989 \$4974 \$4828 \$4985 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7004 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7005 VPWR \$4985 VGND VPWR \$5011 \$4492 \$4974 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$7006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7007 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7008 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7010 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7011 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7012 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7013 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7014 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7016 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7017 VPWR \$5021 VGND VPWR mgmt_gpio_in[15] VGND sky130_fd_sc_hd__clkbuf_1
X$7018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7019 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7020 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7023 VPWR \$953 VGND VPWR sram_ro_data[6] VGND sky130_fd_sc_hd__clkbuf_1
X$7024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7025 VPWR \$896 VGND VPWR \$897 VGND sky130_fd_sc_hd__clkbuf_1
X$7026 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7027 VGND \$897 \$906 \$905 \$918 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7029 VPWR \$906 VGND \$768 VPWR \$935 \$954 \$919 VGND
+ sky130_fd_sc_hd__a31oi_1
X$7030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7031 VGND \$905 \$945 \$954 \$564 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7032 VPWR VGND \$768 VPWR \$935 \$919 \$906 VGND sky130_fd_sc_hd__a21oi_1
X$7033 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7035 VPWR VGND \$720 \$945 \$935 \$955 \$768 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7038 VGND \$877 \$599 \$381 \$811 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$7039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7040 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7041 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7044 VPWR \$898 VGND VPWR \$565 VGND sky130_fd_sc_hd__clkbuf_1
X$7045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7047 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7048 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7049 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7050 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7051 VPWR \$956 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$7052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7056 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7057 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7058 VPWR \$957 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$7059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7062 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7063 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7064 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7067 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7068 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7069 VPWR \$921 \$461 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7070 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7071 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7072 VGND \$856 \$909 \$922 \$908 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7073 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7076 VPWR VGND \$701 \$281 \$909 \$908 \$711 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7077 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7078 VPWR VGND VPWR \$958 \$909 VGND sky130_fd_sc_hd__inv_2
X$7079 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7080 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7081 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7082 VGND \$655 \$959 \$922 \$937 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7085 VPWR VGND \$792 \$281 \$959 \$937 \$793 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7087 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7088 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7090 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7092 VGND \$655 \$939 \$961 \$938 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7094 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7095 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7096 VPWR VGND VPWR \$892 \$911 VGND sky130_fd_sc_hd__inv_2
X$7097 VPWR VGND \$892 \$294 \$939 \$938 \$911 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7099 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7100 VPWR \$924 \$858 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7102 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7103 VPWR VGND \$602 \$293 \$963 \$962 \$674 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7104 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7105 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7107 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7108 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7110 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7112 VPWR VGND VPWR \$912 \$893 VGND sky130_fd_sc_hd__inv_2
X$7113 VPWR VGND \$884 \$925 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$7114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7116 VGND \$655 \$900 \$605 \$926 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$7117 VPWR VGND \$912 \$281 \$900 \$926 \$893 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7118 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7119 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7120 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7122 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7123 VPWR \$928 VGND VPWR \$946 VGND sky130_fd_sc_hd__clkbuf_1
X$7124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7126 VGND \$655 \$1152 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$7127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7128 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7129 VPWR \$913 VGND \$1507 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$7130 VPWR VPWR VGND \$913 \$607 VGND sky130_fd_sc_hd__clkbuf_2
X$7131 VGND \$655 \$947 \$771 \$965 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7135 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7136 VGND \$940 \$964 \$948 \$848 \$347 \$579 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7138 VPWR \$929 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7140 VPWR VGND VPWR \$948 \$730 VGND sky130_fd_sc_hd__inv_2
X$7141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7142 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7143 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7144 VPWR \$929 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7145 VGND \$516 \$949 \$771 \$967 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7146 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7147 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7150 VGND \$516 \$894 \$435 \$901 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7153 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7154 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7155 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7156 VPWR VGND \$713 \$281 \$950 \$969 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$7157 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7160 VPWR VPWR VGND \$966 \$466 VGND sky130_fd_sc_hd__clkbuf_2
X$7161 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7163 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7165 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7166 VPWR \$931 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7168 VGND \$930 \$982 \$931 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7169 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7171 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7172 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7173 VGND \$888 \$970 \$951 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7174 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7176 VGND \$971 \$289 \$1049 \$942 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$7177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7178 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7179 VGND \$516 \$952 \$466 \$972 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7180 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7181 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7187 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7188 VGND \$836 \$974 \$886 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7190 VPWR VGND VPWR \$973 \$322 VGND sky130_fd_sc_hd__inv_2
X$7191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7192 VGND \$677 \$672 \$914 \$973 \$932 VPWR VPWR VGND sky130_fd_sc_hd__a31o_1
X$7193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7194 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7197 VPWR VGND \$903 VPWR \$322 \$745 \$902 VGND sky130_fd_sc_hd__a21o_1
X$7198 VPWR \$777 VGND \$808 \$975 VPWR \$943 VGND sky130_fd_sc_hd__o21ai_2
X$7199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7200 VGND \$976 \$934 \$915 \$933 \$808 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2a_2
X$7201 VGND \$933 \$915 \$943 \$777 \$902 VPWR VPWR VGND sky130_fd_sc_hd__o31a_1
X$7202 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7203 VPWR \$943 VPWR VGND \$934 \$777 \$808 VGND sky130_fd_sc_hd__or3_2
X$7204 VGND \$746 \$915 \$934 \$904 \$889 \$916 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$7205 VPWR VGND VPWR \$915 \$944 VGND sky130_fd_sc_hd__inv_2
X$7206 VPWR \$915 VGND \$934 \$916 VPWR \$904 VGND sky130_fd_sc_hd__o21ai_2
X$7207 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7208 VPWR \$943 \$944 VGND \$759 VPWR \$1012 \$698 VGND sky130_fd_sc_hd__or4_2
X$7209 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7210 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7211 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7214 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7215 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7216 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7217 VPWR VGND \$1039 \$1051 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$7218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7219 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7220 VPWR \$1068 VGND VPWR \$573 \$308 VGND sky130_fd_sc_hd__and2b_1
X$7221 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7222 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7225 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7226 VGND \$1132 \$720 \$955 \$564 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7227 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7228 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7230 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7231 VGND \$1092 \$623 \$999 \$1078 \$1079 \$790 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$7232 VPWR \$1069 VPWR VGND \$720 \$999 VGND sky130_fd_sc_hd__nand2_1
X$7233 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7236 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7237 VPWR \$1052 VGND \$1069 \$623 VPWR VGND sky130_fd_sc_hd__or2_1
X$7238 VPWR VGND \$1052 \$1014 \$1015 \$1040 \$574 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7240 VGND \$1041 \$1014 \$387 \$1040 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$7241 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7244 VPWR VGND VPWR \$1053 \$1055 VGND sky130_fd_sc_hd__inv_2
X$7245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7246 VPWR VGND \$1053 \$1054 \$986 \$1043 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7247 VGND \$565 \$864 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$7248 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7249 VGND \$1054 \$780 \$1000 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7252 VPWR VGND \$1053 \$1056 \$1002 \$978 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7253 VGND \$1056 \$986 \$1057 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7254 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7255 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7256 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7257 VPWR \$986 VPWR \$1057 VGND \$1085 \$1002 VGND sky130_fd_sc_hd__o21a_1
X$7258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7259 VPWR \$1044 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$7260 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7261 VGND \$1070 \$1093 \$1086 \$1016 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7262 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7263 VPWR \$1070 VGND VPWR \$1044 VGND sky130_fd_sc_hd__clkbuf_1
X$7264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7265 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7266 VPWR VGND VPWR \$1072 \$193 VGND sky130_fd_sc_hd__inv_2
X$7267 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7269 VGND \$856 \$1074 \$891 \$1073 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7270 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7271 VPWR VGND \$1087 \$293 \$1074 \$1073 \$1088 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7272 VPWR VGND VPWR \$1087 \$1088 VGND sky130_fd_sc_hd__inv_2
X$7273 VPWR VGND \$1087 \$183 \$1094 \$1095 \$1088 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7275 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7277 VPWR VGND VPWR \$1163 \$1074 VGND sky130_fd_sc_hd__inv_2
X$7278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7279 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7280 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7282 VPWR \$1032 VGND \$1058 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$7283 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7285 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7286 VPWR \$1075 VGND VPWR \$334 \$456 \$1081 \$1058 VGND
+ sky130_fd_sc_hd__o22a_1
X$7287 VPWR \$1081 \$979 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7288 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7289 VPWR \$867 VPWR VGND \$1059 \$1034 \$345 VGND sky130_fd_sc_hd__or3_1
X$7290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7291 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7293 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7294 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7298 VPWR VGND \$980 \$1076 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$7299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7301 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7302 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7303 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7304 VGND \$655 \$981 \$961 \$1006 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7305 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7306 VPWR VGND VPWR \$1097 \$981 VGND sky130_fd_sc_hd__inv_2
X$7307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7309 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7310 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7312 VPWR \$1033 VGND \$1060 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$7313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7315 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7316 VPWR VGND \$1061 \$1030 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$7317 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7318 VPWR \$1077 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7319 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7320 VPWR \$1098 VGND VPWR \$1077 \$1089 \$1028 \$1114 VGND
+ sky130_fd_sc_hd__o22a_1
X$7321 VPWR VGND \$912 \$293 \$1061 \$1021 \$893 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7322 VGND \$1047 \$1098 \$925 \$859 \$686 \$473 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7324 VPWR \$4275 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7327 VPWR \$345 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7328 VPWR \$1046 VPWR VGND \$1034 \$1257 \$345 VGND sky130_fd_sc_hd__or3_1
X$7329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7330 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7331 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7335 VPWR \$910 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7336 VGND \$1082 \$1075 \$910 \$1089 \$755 \$253 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7338 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7341 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7342 VGND \$655 \$1035 \$771 \$1062 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7344 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7347 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7348 VGND \$1067 \$870 \$1090 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7351 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7352 VPWR VGND VPWR \$1701 \$894 VGND sky130_fd_sc_hd__inv_2
X$7353 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7355 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7358 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7359 VPWR \$1063 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7360 VGND \$636 \$894 \$1063 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7363 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7364 VGND \$873 \$1093 \$1064 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7366 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7367 VPWR \$1064 \$950 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7368 VPWR \$1083 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7370 VPWR VGND VPWR \$1563 \$982 VGND sky130_fd_sc_hd__inv_2
X$7371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7374 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7377 VPWR VPWR VGND \$1066 \$246 VGND sky130_fd_sc_hd__clkbuf_2
X$7378 VGND \$667 \$950 \$1036 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7380 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7381 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7384 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7385 VGND \$1026 \$1049 \$1119 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7389 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7391 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7393 VPWR VGND VPWR \$1037 \$1067 VGND sky130_fd_sc_hd__inv_2
X$7394 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7395 VPWR VGND VPWR \$289 \$1038 VGND sky130_fd_sc_hd__inv_4
X$7396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7399 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7400 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7401 VGND \$516 \$895 \$466 \$1084 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$7402 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7405 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7406 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7408 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7409 VGND \$516 \$944 \$246 \$976 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7410 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7411 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7412 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7417 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7420 VPWR \$2319 VGND VPWR sram_ro_data[29] VGND sky130_fd_sc_hd__clkbuf_1
X$7421 VPWR VGND VPWR \$2381 \$2387 VGND sky130_fd_sc_hd__inv_2
X$7422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7424 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7425 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7426 VPWR VGND VPWR \$2407 \$2362 VGND sky130_fd_sc_hd__inv_2
X$7427 VPWR \$2362 VGND \$2154 \$1979 VPWR VGND sky130_fd_sc_hd__or2_1
X$7428 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7430 VGND \$2211 \$2389 \$2408 \$2388 \$2154 \$1897 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$7431 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7432 VPWR \$2187 VGND \$2435 VPWR \$2352 VGND sky130_fd_sc_hd__nor2_1
X$7433 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7434 VGND \$2233 \$2154 \$2363 \$2187 \$2362 \$1897 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_4
X$7435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7436 VPWR \$2409 VGND \$2154 VPWR \$1962 VGND sky130_fd_sc_hd__nor2_1
X$7437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7439 VPWR VGND VPWR \$2336 \$2214 VGND sky130_fd_sc_hd__inv_4
X$7440 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7441 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7442 VPWR \$2364 VGND \$2235 \$2353 VPWR VGND sky130_fd_sc_hd__or2_1
X$7443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7444 VGND \$2410 \$2412 \$2365 \$2425 \$1899 \$2390 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2111o_2
X$7445 VPWR \$2365 VPWR VGND \$2354 \$2311 \$2364 VGND sky130_fd_sc_hd__or3_1
X$7446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7447 VPWR \$2425 VGND \$1933 \$2391 VPWR VGND sky130_fd_sc_hd__or2_1
X$7448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7450 VPWR \$2198 VGND \$2320 VPWR \$2337 VGND sky130_fd_sc_hd__nor2_1
X$7451 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7452 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7453 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7454 VPWR VGND VPWR \$2171 \$2337 VGND sky130_fd_sc_hd__inv_2
X$7455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7456 VPWR \$1981 VGND \$2234 VPWR \$2337 VGND sky130_fd_sc_hd__nor2_1
X$7457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7458 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7459 VPWR \$2443 VGND \$1921 \$2392 VPWR VGND sky130_fd_sc_hd__or2_1
X$7460 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7461 VPWR \$2413 VGND \$1981 \$2393 VPWR VGND sky130_fd_sc_hd__or2_1
X$7462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7463 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7464 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7465 VPWR \$2414 VGND \$2058 \$2394 VPWR VGND sky130_fd_sc_hd__or2_1
X$7466 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7469 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7471 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7472 VPWR VGND \$1771 \$281 \$2338 \$2313 \$1815 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7476 VPWR VGND VPWR \$2382 \$2338 VGND sky130_fd_sc_hd__inv_2
X$7477 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7478 VGND \$2395 \$2381 \$1556 \$686 \$921 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$7479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7481 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7483 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7484 VPWR VGND VPWR \$2321 \$2322 VGND sky130_fd_sc_hd__inv_2
X$7485 VGND \$856 \$2339 \$1861 \$2340 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7488 VPWR VPWR VGND \$2396 \$2322 VGND sky130_fd_sc_hd__clkbuf_2
X$7489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7490 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7491 VPWR \$2396 VGND \$2355 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$7492 VPWR VGND VPWR \$2298 \$2339 VGND sky130_fd_sc_hd__inv_2
X$7493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7494 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7495 VPWR \$1570 VGND VPWR \$2366 \$1401 VGND sky130_fd_sc_hd__or2_4
X$7496 VPWR \$1598 VGND VPWR \$2372 \$1401 VGND sky130_fd_sc_hd__or2_4
X$7497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7499 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7500 VPWR \$1598 VGND VPWR \$2355 \$1356 VGND sky130_fd_sc_hd__or2_4
X$7501 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7502 VPWR \$2356 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7503 VPWR \$1598 VGND VPWR \$2384 \$1257 VGND sky130_fd_sc_hd__or2_4
X$7504 VGND \$2367 \$2356 \$769 \$1058 \$1556 \$2310 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7506 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7507 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7511 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7512 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7513 VGND \$2370 \$2343 \$725 \$2369 \$2357 \$2296 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7514 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7515 VGND \$2371 \$2344 \$601 \$2369 \$2357 \$2122 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7516 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7517 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7518 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7519 VGND \$2368 \$2088 \$2355 \$1116 \$1236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$7520 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7521 VGND \$2359 \$1763 \$2341 \$3042 \$2355 \$2298 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7524 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7526 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7530 VPWR \$2373 VGND VPWR \$1419 \$1643 \$2323 \$2372 VGND
+ sky130_fd_sc_hd__o22a_1
X$7531 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7532 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7534 VGND \$2398 \$2373 \$2297 \$2384 \$1625 \$2397 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7535 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7536 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7538 VGND \$1733 \$2359 \$2285 \$2113 \$2325 \$2360 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7541 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7542 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7543 VPWR VGND VPWR \$1698 \$2317 \$2398 \$2385 \$2361 VGND
+ sky130_fd_sc_hd__and4_1
X$7544 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7545 VPWR \$2361 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7546 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7547 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7548 VGND \$2385 \$1234 \$576 \$379 \$2386 \$2400 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7549 VGND \$2374 \$560 \$534 \$2375 \$2615 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2a_2
X$7550 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7552 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7553 VPWR \$2399 VGND VPWR \$2324 \$1956 \$1943 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$7554 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7555 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7559 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7561 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7565 VPWR \$2347 VPWR VGND \$1128 \$1882 \$1679 VGND sky130_fd_sc_hd__or3_1
X$7566 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7567 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7568 VGND \$2347 \$2316 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7569 VPWR \$2417 VPWR VGND \$1128 \$1384 \$1705 VGND sky130_fd_sc_hd__or3_1
X$7570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7571 VGND \$2349 \$2724 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7572 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7573 VPWR \$1448 \$2418 \$1415 VPWR VGND \$1384 \$1705 VGND
+ sky130_fd_sc_hd__or4_1
X$7574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7575 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7576 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7578 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7579 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7580 VPWR \$2376 VGND \$2277 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$7581 VPWR \$2331 VGND \$2277 \$1780 VPWR VGND sky130_fd_sc_hd__or2_1
X$7582 VGND \$2376 \$2809 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7583 VPWR \$2332 VGND \$1782 \$2231 VPWR VGND sky130_fd_sc_hd__or2_1
X$7584 VPWR \$2290 VGND \$2231 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$7585 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7587 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7588 VGND \$1152 \$2378 \$2255 \$2377 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7589 VPWR VGND \$2401 \$1179 \$2378 \$2377 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7590 VPWR VGND VPWR \$2360 \$2378 VGND sky130_fd_sc_hd__inv_2
X$7591 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7594 VPWR VGND VPWR \$2401 \$2334 VGND sky130_fd_sc_hd__inv_2
X$7595 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7600 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7601 VPWR VGND \$2402 \$2403 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$7602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7603 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7605 VPWR \$2848 \$2350 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7606 VPWR VGND \$2127 \$1171 \$2404 \$2420 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7608 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7611 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7612 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7613 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7614 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7615 VPWR VGND \$2127 \$386 \$2379 \$2380 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7616 VGND \$1152 \$2379 \$2232 \$2380 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7617 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7618 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7619 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7621 VPWR \$2421 VGND VPWR \$2405 VGND sky130_fd_sc_hd__clkbuf_1
X$7622 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7623 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7629 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7630 VPWR VGND VPWR \$1964 \$1959 VGND sky130_fd_sc_hd__inv_2
X$7631 VPWR \$1959 VGND VPWR sram_ro_data[23] VGND sky130_fd_sc_hd__clkbuf_1
X$7632 VGND \$1973 \$1945 \$1974 \$1514 \$1473 VPWR VPWR VGND
+ sky130_fd_sc_hd__a22o_2
X$7633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7634 VGND \$1930 \$1945 \$1376 \$1974 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$7635 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7636 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7638 VPWR \$1896 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$7639 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7640 VPWR \$1930 VGND VPWR \$1896 VGND sky130_fd_sc_hd__clkbuf_1
X$7641 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7642 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7643 VPWR \$1975 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7644 VGND \$1976 \$1975 \$1945 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7645 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7647 VPWR \$1933 VGND \$1960 VPWR \$1962 VGND sky130_fd_sc_hd__nor2_1
X$7648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7649 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7650 VPWR VGND \$1960 VPWR \$1961 VGND sky130_fd_sc_hd__clkbuf_4
X$7651 VPWR \$1918 VGND \$1931 \$1932 \$2024 VPWR \$1919 VGND
+ sky130_fd_sc_hd__nor4_1
X$7652 VPWR \$1898 VPWR VGND \$2236 \$1933 \$1899 VGND sky130_fd_sc_hd__or3_1
X$7653 VPWR \$1932 VGND \$1960 VPWR \$1963 VGND sky130_fd_sc_hd__nor2_1
X$7654 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7655 VGND \$1977 \$1978 \$2025 \$1886 \$1918 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$7656 VPWR \$1918 VGND \$1920 VPWR \$1897 VGND sky130_fd_sc_hd__nor2_1
X$7657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7658 VPWR \$1946 VGND \$1920 \$1963 VPWR VGND sky130_fd_sc_hd__or2_1
X$7659 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7660 VPWR \$1980 VGND \$1920 \$1979 VPWR VGND sky130_fd_sc_hd__or2_1
X$7661 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7662 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7664 VPWR VGND VPWR \$1886 \$1980 VGND sky130_fd_sc_hd__inv_2
X$7665 VPWR \$1921 VGND \$1920 VPWR \$1962 VGND sky130_fd_sc_hd__nor2_1
X$7666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7667 VPWR \$1934 VGND \$1921 \$1901 VPWR VGND sky130_fd_sc_hd__or2_1
X$7668 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7669 VPWR \$1982 VGND \$1981 \$1934 VPWR VGND sky130_fd_sc_hd__or2_1
X$7670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7671 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7673 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7674 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7676 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7677 VPWR VGND \$1725 \$1398 \$1922 \$1935 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7678 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7679 VGND \$856 \$1903 \$1750 \$1936 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7681 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7682 VPWR VPWR VGND \$1902 \$387 VGND sky130_fd_sc_hd__clkbuf_2
X$7683 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7684 VPWR VGND \$1923 \$200 \$1903 \$1936 \$1924 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7686 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7687 VPWR VGND \$1923 \$281 \$1983 \$2003 \$1924 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7688 VPWR \$1852 \$1903 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7689 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7690 VPWR VPWR VGND \$1984 \$1924 VGND sky130_fd_sc_hd__clkbuf_2
X$7691 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7692 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7693 VPWR \$1984 VGND \$1729 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$7694 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7696 VGND \$856 \$1905 \$1370 \$1904 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7697 VPWR \$1947 VGND VPWR \$1964 \$1554 \$1451 \$1297 VGND
+ sky130_fd_sc_hd__o22a_1
X$7698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7699 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7701 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7702 VPWR \$1948 \$1905 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7705 VGND \$1906 \$927 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$7706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7707 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7710 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7711 VGND \$463 \$1863 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$7712 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7713 VPWR \$1925 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7714 VPWR \$1937 VGND VPWR \$778 \$1114 \$1925 \$1219 VGND
+ sky130_fd_sc_hd__o22a_1
X$7715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7716 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7717 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7719 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7720 VPWR \$1949 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7721 VGND \$1836 \$1937 \$1949 \$1466 \$1556 \$2166 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7724 VGND \$1938 \$1864 \$1907 \$1715 \$1754 \$1097 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7726 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7727 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7729 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7730 VPWR \$1985 VGND VPWR \$1965 \$1966 \$1851 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$7731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7732 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7733 VPWR \$1986 VGND VPWR \$1852 \$1967 \$1851 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$7734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7736 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7740 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7741 VPWR \$3163 VGND VPWR \$1907 \$1613 \$1427 \$1421 VGND
+ sky130_fd_sc_hd__o22a_1
X$7742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7744 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7745 VPWR \$1952 VGND VPWR \$616 \$2045 \$1968 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$7746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7750 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7751 VPWR \$1988 VGND VPWR \$1427 \$1956 \$1869 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$7752 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7753 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7754 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7755 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7757 VPWR \$345 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7758 VPWR \$1911 VGND \$1890 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$7759 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7760 VPWR VGND VPWR \$1989 \$1910 VGND sky130_fd_sc_hd__inv_2
X$7761 VGND \$1152 \$1910 \$1627 \$1926 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7763 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7765 VPWR \$1990 VGND VPWR \$1927 \$1879 \$645 \$347 VGND
+ sky130_fd_sc_hd__o22a_1
X$7766 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7767 VGND \$1152 \$1991 \$1627 \$1969 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$7768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7769 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7770 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7773 VGND \$1844 \$1928 \$1883 \$1870 \$1912 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$7774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7775 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7776 VPWR \$1940 VGND VPWR \$554 \$1562 \$1869 \$1890 VGND
+ sky130_fd_sc_hd__o22a_1
X$7777 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7780 VPWR \$1992 VPWR VGND \$1449 \$1882 \$1679 VGND sky130_fd_sc_hd__or3_1
X$7781 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7782 VGND \$1992 \$1967 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7783 VPWR \$1941 VPWR VGND \$1384 \$1449 \$1679 VGND sky130_fd_sc_hd__or3_1
X$7784 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7785 VPWR \$1448 \$1970 \$1415 VPWR VGND \$1882 \$1705 VGND
+ sky130_fd_sc_hd__or4_1
X$7786 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7787 VGND \$1970 \$1987 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7788 VPWR \$1942 VPWR VGND \$1384 \$1449 \$1705 VGND sky130_fd_sc_hd__or3_1
X$7789 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7790 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7791 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7792 VPWR \$1993 VPWR VGND \$1797 \$1746 \$1782 VGND sky130_fd_sc_hd__or3_1
X$7793 VGND \$1913 \$2005 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7794 VGND \$1971 \$2047 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7795 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7796 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7797 VPWR \$1662 \$2081 \$1308 VPWR VGND \$1814 \$1782 VGND
+ sky130_fd_sc_hd__or4_1
X$7798 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7799 VPWR \$1662 \$1944 \$1308 VPWR VGND \$1746 \$1766 VGND
+ sky130_fd_sc_hd__or4_1
X$7800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7801 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7802 VPWR \$1662 \$1994 \$1308 VPWR VGND \$1746 \$1782 VGND
+ sky130_fd_sc_hd__or4_1
X$7803 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7805 VPWR \$1782 VGND VPWR \$2007 \$1533 VGND sky130_fd_sc_hd__or2_4
X$7806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7808 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7809 VPWR \$1929 VGND \$1766 \$1533 VPWR VGND sky130_fd_sc_hd__or2_1
X$7810 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7811 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7812 VGND \$1929 \$1536 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7813 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7815 VPWR VGND VPWR \$1915 \$1857 VGND sky130_fd_sc_hd__inv_2
X$7816 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7817 VPWR \$1943 \$1858 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7820 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7822 VGND \$1335 \$927 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$7823 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7824 VPWR \$1995 VGND \$2117 \$927 VPWR VGND sky130_fd_sc_hd__or2_1
X$7825 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7828 VGND \$516 \$1996 \$1273 \$1958 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7829 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7830 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7831 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7832 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7834 VGND \$516 \$1895 \$1273 \$1916 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$7835 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7836 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7837 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7838 VPWR mgmt_gpio_in[5] VPWR VGND \$1997 VGND sky130_fd_sc_hd__buf_4
X$7839 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7843 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7844 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7845 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7846 VPWR \$1655 \$2038 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7847 VPWR \$2013 \$2012 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7848 VPWR VGND \$1514 \$2056 \$2040 \$2039 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7850 VGND \$2056 \$2057 \$1860 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7852 VGND \$1973 \$2221 \$2040 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$7853 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7854 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7855 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7857 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7858 VPWR \$2024 \$2014 VPWR \$2001 \$1999 \$1960 VGND \$1897 VGND
+ sky130_fd_sc_hd__o221ai_1
X$7859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7860 VPWR \$1961 VGND \$1999 \$2015 VPWR VGND sky130_fd_sc_hd__or2_1
X$7861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7862 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7863 VPWR VGND \$1998 VPWR \$1919 \$1960 VGND sky130_fd_sc_hd__nor2_2
X$7864 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7866 VPWR \$2025 VGND \$1899 \$1932 VPWR VGND sky130_fd_sc_hd__or2_1
X$7867 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7868 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7870 VGND \$2000 \$1946 \$2016 \$1931 \$2002 \$2001 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$7871 VPWR \$2016 VGND \$1920 \$1998 VPWR VGND sky130_fd_sc_hd__or2_1
X$7872 VPWR VGND VPWR \$2041 \$2016 VGND sky130_fd_sc_hd__inv_2
X$7873 VPWR \$1920 VGND \$2002 \$2015 VPWR VGND sky130_fd_sc_hd__or2_1
X$7874 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7875 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7876 VPWR VGND VPWR \$2017 \$1946 VGND sky130_fd_sc_hd__inv_2
X$7877 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7878 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7879 VPWR VPWR \$1897 VGND \$2026 \$2027 \$2000 VGND sky130_fd_sc_hd__o21ai_1
X$7880 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7881 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7882 VPWR \$2058 VGND \$2026 VPWR \$1979 VGND sky130_fd_sc_hd__nor2_1
X$7883 VPWR \$2059 VGND \$2058 \$1982 VPWR VGND sky130_fd_sc_hd__or2_1
X$7884 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7886 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7887 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7888 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7889 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7890 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7892 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7893 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7894 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7895 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7896 VPWR VGND VPWR \$1923 \$1924 VGND sky130_fd_sc_hd__inv_2
X$7897 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7898 VGND \$856 \$1983 \$1370 \$2003 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$7899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7901 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7903 VPWR \$2018 \$1983 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$7904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7907 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7908 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7911 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7912 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7914 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7915 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7920 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7921 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7929 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7930 VGND \$2061 \$1985 \$2060 \$2043 \$1914 \$631 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7931 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7932 VPWR \$2029 VGND VPWR \$1989 \$1890 \$631 \$1060 VGND
+ sky130_fd_sc_hd__o22a_1
X$7933 VPWR \$1490 VGND VPWR \$2113 \$1435 VGND sky130_fd_sc_hd__or2_4
X$7934 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7935 VPWR \$2028 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$7936 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7937 VGND \$2030 \$631 \$2005 \$2028 \$2019 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$7938 VGND \$2062 \$2063 \$2030 \$2044 VPWR \$580 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$7939 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7940 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7941 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7942 VGND \$2019 \$1986 \$703 \$1953 \$1987 \$1202 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7943 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7944 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7945 VPWR \$2006 VGND VPWR \$2018 \$1967 \$1948 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$7946 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7947 VGND \$2032 \$2006 \$616 \$1953 \$1987 \$1427 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7948 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7949 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7950 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$7951 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$7952 VGND \$2064 \$2078 \$2077 \$2034 VPWR \$519 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$7953 VGND \$1841 \$2004 \$1968 \$1558 \$1867 \$2033 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7954 VGND \$2034 \$1909 \$2020 \$2065 \$2046 \$1968 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7955 VGND \$1988 \$2020 \$2047 \$2048 \$661 \$2042 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$7956 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7957 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7958 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7959 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7960 VGND \$2044 \$2035 \$2066 \$2065 \$2046 \$1529 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$7961 VPWR \$2021 VGND VPWR \$1202 \$1956 \$1989 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$7962 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7963 VPWR \$2035 VGND VPWR \$1611 \$1793 \$1989 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$7964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7965 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7966 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7970 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7971 VPWR VGND \$2049 \$200 \$1991 \$1969 \$2050 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7972 VPWR VGND VPWR \$2066 \$1991 VGND sky130_fd_sc_hd__inv_2
X$7973 VPWR VGND \$2049 \$281 \$2051 \$2067 \$2050 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$7974 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7975 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7976 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$7978 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7979 VPWR VGND VPWR \$2020 \$2051 VGND sky130_fd_sc_hd__inv_2
X$7980 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$7982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7983 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7984 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7985 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$7986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7987 VGND \$2036 \$1939 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7988 VPWR \$2036 VPWR VGND \$1128 \$1384 \$1679 VGND sky130_fd_sc_hd__or3_1
X$7989 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$7990 VGND \$1941 \$1953 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7991 VGND \$2079 \$2065 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7992 VGND \$1942 \$2046 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$7993 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$7994 VPWR \$1662 \$2052 \$1308 VPWR VGND \$1814 \$1766 VGND
+ sky130_fd_sc_hd__or4_1
X$7995 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$7996 VPWR \$2037 VPWR VGND \$1663 \$1746 \$1782 VGND sky130_fd_sc_hd__or3_1
X$7997 VGND \$2037 \$2096 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$7998 VGND \$1993 \$2048 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$7999 VPWR \$1662 \$2126 \$1308 VPWR VGND \$1783 \$1780 VGND
+ sky130_fd_sc_hd__or4_1
X$8000 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8001 VGND \$1944 \$1951 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$8002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8003 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8004 VPWR \$1783 \$1308 VGND \$1662 VPWR \$2483 \$1766 VGND
+ sky130_fd_sc_hd__or4_2
X$8005 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8006 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8007 VGND \$2022 \$1956 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$8008 VGND \$2054 \$880 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$8009 VPWR \$2008 VGND \$2180 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$8010 VPWR \$2022 VGND \$1782 \$1801 VPWR VGND sky130_fd_sc_hd__or2_1
X$8011 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8013 VPWR VGND \$1681 VPWR \$2008 VGND sky130_fd_sc_hd__clkbuf_4
X$8014 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8015 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8016 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8018 VPWR VGND \$1680 \$354 \$2009 \$2010 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8019 VPWR \$2053 \$2009 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8021 VGND \$516 \$2009 \$1273 \$2010 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8022 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8023 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8025 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8027 VPWR VGND \$1310 VPWR \$1995 VGND sky130_fd_sc_hd__clkbuf_4
X$8028 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8029 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8030 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8031 VPWR VGND \$1311 \$184 \$1996 \$1958 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8032 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8033 VGND \$2055 \$184 \$1996 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$8034 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8035 VGND \$516 \$2068 \$1273 \$2023 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8036 VPWR \$2023 VGND VPWR \$2055 \$1363 \$2068 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$8037 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8038 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8041 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8042 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8045 VPWR VGND wb_dat_o[26] VPWR \$5189 VGND sky130_fd_sc_hd__buf_2
X$8046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8047 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8048 VGND \$4907 \$4651 \$5199 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$8049 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8050 VPWR \$5199 VGND VPWR \$4907 \$5076 \$2057 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$8051 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8052 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8054 VPWR VGND \$4509 VPWR \$5218 VGND sky130_fd_sc_hd__clkbuf_4
X$8055 VPWR \$4930 \$5180 \$4917 VPWR VGND \$4941 \$5147 VGND
+ sky130_fd_sc_hd__or4_1
X$8056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8057 VGND \$5180 \$1897 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$8058 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8059 VGND \$4853 \$4698 \$4891 \$4881 \$4864 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$8060 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8062 VPWR \$5181 VGND \$5190 \$4863 VPWR VGND sky130_fd_sc_hd__or2_1
X$8063 VPWR VGND VPWR \$5169 \$5190 VGND sky130_fd_sc_hd__inv_2
X$8064 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8065 VPWR \$5169 VGND \$5170 \$5110 VPWR \$4854 VGND sky130_fd_sc_hd__o21ai_2
X$8066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8067 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8068 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8069 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8070 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8071 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8072 VPWR \$3857 \$2571 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8073 VGND \$5200 \$5219 \$2390 \$5220 \$5201 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$8074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8075 VGND \$5233 \$5220 \$5219 \$3857 \$5200 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$8076 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8077 VPWR \$5361 VGND \$4772 \$4855 VPWR VGND sky130_fd_sc_hd__or2_1
X$8078 VPWR \$5222 VGND \$5221 \$4772 VPWR VGND sky130_fd_sc_hd__or2_1
X$8079 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8080 VPWR \$5191 VGND \$5222 \$5113 VPWR VGND sky130_fd_sc_hd__or2_1
X$8081 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8082 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8083 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8084 VPWR \$5182 VPWR VGND \$5106 \$3663 \$5191 VGND sky130_fd_sc_hd__or3_1
X$8085 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8086 VPWR \$3411 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8087 VPWR \$4777 VGND \$5213 \$5336 \$3117 VPWR \$3411 VGND
+ sky130_fd_sc_hd__nor4_1
X$8088 VPWR \$5201 VGND \$5182 \$4153 VPWR VGND sky130_fd_sc_hd__or2_1
X$8089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8090 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8091 VPWR VPWR VGND \$4715 \$5002 VGND sky130_fd_sc_hd__clkbuf_2
X$8092 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8094 VPWR \$5234 VPWR VGND \$5183 \$5202 \$5223 VGND sky130_fd_sc_hd__or3_1
X$8095 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8096 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8099 VPWR \$4520 VPWR VGND \$4676 \$4758 VGND sky130_fd_sc_hd__or2_2
X$8100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8102 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8103 VPWR \$5214 VPWR VGND \$5203 \$5235 VGND sky130_fd_sc_hd__or2_2
X$8104 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8105 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8106 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8107 VPWR \$5218 VGND \$5235 \$5224 VPWR VGND sky130_fd_sc_hd__or2_1
X$8108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8110 VPWR \$5236 VGND \$5225 \$5116 VPWR VGND sky130_fd_sc_hd__or2_1
X$8111 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8112 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8113 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8114 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8115 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8117 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8118 VPWR \$5215 \$5204 VGND \$5226 VPWR \$4934 \$5176 VGND
+ sky130_fd_sc_hd__or4_2
X$8119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8120 VPWR VGND VPWR \$5203 \$5204 VGND sky130_fd_sc_hd__inv_2
X$8121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8123 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8124 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8125 VGND \$2777 \$5185 \$4811 \$5205 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$8126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8127 VPWR VGND \$5192 \$4774 \$5185 \$5205 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8130 VPWR VGND \$5185 \$3312 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8131 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8132 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8135 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8136 VPWR \$3734 \$5227 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8138 VPWR VGND \$5097 \$184 \$5228 \$5237 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8141 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8142 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8143 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8146 VPWR \$5238 VGND \$1125 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$8147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8149 VGND \$4761 \$5193 \$4994 \$5206 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8150 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8151 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8154 VPWR \$5186 VGND \$1089 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$8155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8156 VPWR VGND \$5193 \$2917 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8157 VPWR VGND \$5229 \$354 \$5217 \$5216 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8158 VPWR VGND \$5207 VPWR \$5186 VGND sky130_fd_sc_hd__clkbuf_4
X$8159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8162 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8163 VPWR \$5239 VGND \$1625 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$8164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8167 VPWR \$5240 VGND \$2162 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$8168 VPWR \$4294 \$5217 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8169 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8170 VPWR VGND \$5230 \$2498 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8171 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8172 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8174 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8175 VPWR VGND \$5044 \$1594 \$5231 \$5241 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8176 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8178 VPWR VGND VPWR \$3004 \$5231 VGND sky130_fd_sc_hd__inv_2
X$8179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8182 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8183 VGND \$4761 \$5194 \$4850 \$5208 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8184 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8185 VPWR VGND \$5194 \$2163 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8189 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8190 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8192 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8193 VPWR VGND VPWR \$5228 \$1099 VGND sky130_fd_sc_hd__inv_4
X$8194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8195 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8197 VPWR \$4293 \$5254 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8200 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8201 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8204 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8205 VGND \$4764 \$5195 \$5006 \$5209 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8207 VPWR \$4088 \$5255 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8208 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8209 VPWR \$4030 \$5195 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8210 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8211 VPWR VGND \$5044 \$184 \$5195 \$5209 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8212 VGND \$4764 \$5187 \$5006 \$5210 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$8213 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8214 VPWR VGND \$5044 \$542 \$5187 \$5210 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8216 VPWR \$2862 \$5187 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$8217 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8218 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8220 VPWR VGND VPWR \$3899 \$5196 VGND sky130_fd_sc_hd__inv_2
X$8221 VGND \$4764 \$5196 \$5006 \$5197 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$8222 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8223 VPWR VGND \$5046 \$4774 \$5196 \$5197 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8225 VGND \$4764 \$5198 \$5006 \$5232 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$8226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8227 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8228 VPWR VGND \$5198 \$3162 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8229 VPWR \$5046 \$4998 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8230 VGND \$4764 \$5177 \$4828 \$5173 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$8231 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8233 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8234 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8235 VPWR \$3611 \$4239 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$8236 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8237 VGND \$4764 \$5161 \$5298 \$5188 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8240 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8247 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8249 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8250 VPWR \$5178 VGND VPWR mgmt_gpio_in[16] VGND sky130_fd_sc_hd__clkbuf_1
X$8251 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8255 VGND \$5075 \$5002 \$5564 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$8256 VPWR VGND spimemio_flash_io1_di VPWR \$1091 VGND sky130_fd_sc_hd__buf_2
X$8257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8258 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8259 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8260 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8261 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8262 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8263 VPWR \$5582 VGND VPWR \$5243 \$5439 \$5448 \$2057 VGND
+ sky130_fd_sc_hd__o22a_1
X$8264 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8265 VPWR \$226 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8266 VGND \$5243 \$4651 \$5582 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$8267 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8268 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8269 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8273 VPWR \$5606 VGND \$5509 VPWR \$5147 VGND sky130_fd_sc_hd__nor2_1
X$8274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8275 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8276 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8278 VGND \$5607 \$4061 \$5597 VPWR VPWR VGND sky130_fd_sc_hd__nand2_4
X$8279 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8280 VPWR \$5597 VGND VPWR \$4050 \$4853 VGND sky130_fd_sc_hd__or2_4
X$8281 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8282 VGND \$4757 \$5583 \$5573 \$4078 \$5471 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4bb_4
X$8283 VPWR \$5584 VGND \$5471 \$5583 VPWR VGND sky130_fd_sc_hd__or2_1
X$8284 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8285 VPWR \$5584 VGND VPWR \$4151 \$5573 VGND sky130_fd_sc_hd__or2_4
X$8286 VPWR \$5574 VGND \$5584 \$5618 VPWR VGND sky130_fd_sc_hd__or2_1
X$8287 VGND \$5574 \$4214 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$8288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8289 VPWR \$5598 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$8290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8292 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8293 VPWR \$5608 VGND VPWR \$5598 VGND sky130_fd_sc_hd__clkbuf_1
X$8294 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8295 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8296 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8298 VPWR VGND \$5504 \$5609 \$5537 \$5555 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8301 VGND \$3711 \$5537 \$1369 \$5610 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$8302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8303 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8305 VPWR VGND \$5504 \$5450 \$5575 \$5639 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8306 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8307 VPWR VGND \$5504 \$5575 \$5485 \$5556 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8308 VPWR \$5599 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$8309 VPWR \$5611 VGND VPWR \$5599 VGND sky130_fd_sc_hd__clkbuf_1
X$8310 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8311 VPWR \$5565 VGND VPWR \$5544 VGND sky130_fd_sc_hd__clkbuf_1
X$8312 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8314 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8315 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8318 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8322 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8324 VPWR \$5149 \$5585 \$5558 \$5586 VGND \$5270 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$8325 VPWR \$5600 \$5612 \$5592 VPWR VGND \$5585 \$1725 VGND
+ sky130_fd_sc_hd__or4_1
X$8326 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8327 VPWR VGND \$5551 VPWR \$5612 VGND sky130_fd_sc_hd__clkbuf_4
X$8328 VPWR VGND VPWR \$5532 \$5423 VGND sky130_fd_sc_hd__inv_2
X$8329 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8330 VPWR VGND \$5613 VPWR \$5614 \$5600 \$5532 VGND sky130_fd_sc_hd__a21oi_1
X$8331 VPWR VGND VPWR \$5339 \$5079 VGND sky130_fd_sc_hd__inv_2
X$8332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8334 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8335 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8337 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8338 VPWR VGND \$5192 \$3732 \$5576 \$5593 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8339 VGND \$2777 \$5576 \$5165 \$5593 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8340 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8341 VPWR VGND VPWR \$5576 \$3444 VGND sky130_fd_sc_hd__inv_4
X$8342 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8344 VPWR VGND \$5559 \$4023 \$5568 \$5587 \$5553 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8345 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8346 VGND \$2777 \$5568 \$5408 \$5587 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8347 VGND \$2777 \$5570 \$5408 \$5569 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8348 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8349 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8351 VPWR VGND \$5568 \$2664 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8352 VPWR VGND VPWR \$5570 \$2685 VGND sky130_fd_sc_hd__inv_4
X$8353 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8354 VGND \$2777 \$5577 \$5408 \$5594 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8355 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8356 VPWR VGND \$5388 \$354 \$5577 \$5594 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8358 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8359 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8361 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8362 VPWR VGND \$5577 \$3675 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$8363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8365 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8367 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8368 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8370 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8372 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8373 VPWR VGND \$5525 \$354 \$5540 \$5560 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8376 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8378 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8379 VPWR VGND \$5498 \$4774 \$5602 \$5615 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8380 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8381 VPWR VGND VPWR \$3723 \$5601 VGND sky130_fd_sc_hd__inv_2
X$8382 VPWR VGND VPWR \$3967 \$5602 VGND sky130_fd_sc_hd__inv_2
X$8383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8384 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8385 VGND \$4761 \$5561 \$5367 \$5571 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$8386 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8387 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8388 VGND \$3952 \$5367 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$8389 VPWR VGND \$5498 \$411 \$5541 \$5588 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8391 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8392 VGND \$4761 \$5541 \$5369 \$5588 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8394 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8395 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8396 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8397 VPWR VGND \$5562 \$184 \$5578 \$5603 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8399 VGND \$4761 \$5578 \$5369 \$5603 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8401 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8402 VPWR \$4628 \$5578 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8405 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8406 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8409 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8410 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8413 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8416 VPWR VGND \$5589 VPWR \$5265 VGND sky130_fd_sc_hd__clkbuf_4
X$8417 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8418 VPWR VGND \$5627 \$354 \$5579 \$5596 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8419 VGND \$4764 \$5579 \$5334 \$5596 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8420 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8421 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8422 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8425 VPWR \$5345 \$5323 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8426 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8427 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8428 VGND \$5515 \$4584 mgmt_gpio_out[32] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$8429 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8430 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8432 VGND \$4764 \$5617 \$5298 \$5580 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8433 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8434 VPWR VGND \$5335 \$411 \$5617 \$5580 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8435 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8436 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8437 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8438 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8439 VPWR VGND \$5335 \$3711 \$5542 \$5563 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8440 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8441 VPWR \$5554 VGND VPWR \$5550 \$4724 \$5572 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$8442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8443 VGND \$5572 \$2908 mgmt_gpio_out[18] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$8444 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8445 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8446 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8448 VPWR VGND \$4483 VPWR mgmt_gpio_in[18] VGND sky130_fd_sc_hd__buf_2
X$8449 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8450 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8451 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8453 VPWR \$1711 VGND VPWR sram_ro_data[21] VGND sky130_fd_sc_hd__clkbuf_1
X$8454 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8455 VPWR VGND VPWR \$1805 \$1131 VGND sky130_fd_sc_hd__inv_2
X$8456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8457 VPWR \$1828 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$8458 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8459 VPWR \$1829 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8461 VGND \$1806 \$1829 \$1684 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$8462 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8464 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8466 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8467 VGND \$1786 \$1769 \$1768 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$8468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8469 VPWR VGND \$1514 \$1976 \$1770 \$1749 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8470 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8471 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8472 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8473 VPWR \$1770 \$1768 VGND VPWR VGND sky130_fd_sc_hd__clkdlybuf4s25_1
X$8474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8476 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8477 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8479 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8481 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8484 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8485 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8486 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8488 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8489 VPWR VGND \$1771 \$293 \$1772 \$1751 \$1815 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8490 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8491 VPWR \$1771 \$1815 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8492 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8495 VGND \$856 \$1833 \$1750 \$1787 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8496 VPWR VGND \$1771 \$183 \$1833 \$1787 \$1815 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8498 VPWR VGND VPWR \$988 \$1772 VGND sky130_fd_sc_hd__inv_2
X$8499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8500 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8501 VGND \$856 \$1773 \$1370 \$1788 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$8502 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8503 VPWR \$1807 \$1540 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8504 VPWR VGND VPWR \$1831 \$1833 VGND sky130_fd_sc_hd__inv_2
X$8505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8507 VPWR VGND VPWR \$1752 \$1774 VGND sky130_fd_sc_hd__inv_2
X$8508 VPWR VGND \$1752 \$200 \$1773 \$1788 \$1774 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8511 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8513 VPWR \$1775 VGND \$1713 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$8514 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8515 VPWR VPWR VGND \$1775 \$1774 VGND sky130_fd_sc_hd__clkbuf_2
X$8516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8519 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8520 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8521 VPWR VGND \$1567 \$281 \$1835 \$1834 \$1568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8526 VPWR VGND VPWR \$1809 \$1836 \$1816 \$1327 \$1808 VGND
+ sky130_fd_sc_hd__and4_1
X$8527 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8530 VGND \$1808 \$336 \$1064 \$848 \$1810 \$1817 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8534 VPWR \$1789 VGND VPWR \$1443 \$1776 \$1115 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$8535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8536 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8539 VPWR \$1837 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8540 VPWR \$1818 VGND VPWR \$638 \$1114 \$1837 \$1810 VGND
+ sky130_fd_sc_hd__o22a_1
X$8541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8542 VPWR \$1283 VGND VPWR \$1819 \$1342 VGND sky130_fd_sc_hd__or2_4
X$8543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8546 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8549 VGND \$1756 \$1818 \$1383 \$1300 \$1819 \$1838 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8550 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8551 VPWR \$1755 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8554 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8555 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8556 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8558 VGND \$1840 \$1117 \$1842 \$1809 \$1791 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$8559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8560 VPWR VGND VPWR \$1791 \$1382 \$1251 \$1777 \$1790 VGND
+ sky130_fd_sc_hd__and4_1
X$8561 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8563 VPWR \$1843 VGND VPWR \$1443 \$1793 \$1820 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$8564 VPWR \$1792 VGND VPWR \$1637 \$1793 \$1778 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$8565 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8566 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8567 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8568 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8569 VGND \$1152 \$1757 \$1627 \$1794 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8570 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8571 VPWR \$1820 \$1757 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8572 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8573 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8576 VGND \$1152 \$1796 \$1627 \$1795 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8577 VPWR VGND \$1572 \$281 \$1796 \$1795 \$1592 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8578 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8579 VPWR \$1846 VGND VPWR \$1821 \$1845 \$215 \$433 VGND
+ sky130_fd_sc_hd__o22a_1
X$8580 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8581 VGND \$1334 \$1812 \$1819 \$320 \$284 \$1847 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$8582 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8583 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8584 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8585 VPWR \$1822 VGND VPWR \$1823 \$1867 \$496 \$320 VGND
+ sky130_fd_sc_hd__o22a_1
X$8586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8590 VPWR VPWR VGND \$1468 \$1066 VGND sky130_fd_sc_hd__clkbuf_2
X$8591 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8593 VPWR \$1824 VGND \$1813 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$8594 VPWR \$1781 VGND \$1779 \$1780 VPWR VGND sky130_fd_sc_hd__or2_1
X$8595 VGND \$1781 \$1715 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$8596 VGND \$1824 \$1754 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$8597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8598 VGND \$1735 \$1793 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$8599 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8600 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8601 VPWR \$1758 VPWR VGND \$1797 \$1746 \$1766 VGND sky130_fd_sc_hd__or3_1
X$8602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8603 VGND \$1825 \$2045 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$8604 VPWR \$1799 VPWR VGND \$1798 \$1746 \$1782 VGND sky130_fd_sc_hd__or3_1
X$8605 VPWR \$1813 VGND \$1783 \$1798 VPWR VGND sky130_fd_sc_hd__or2_1
X$8606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8607 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8608 VPWR \$2080 VPWR VGND \$1574 \$1673 \$1797 VGND sky130_fd_sc_hd__or3_1
X$8609 VPWR \$1574 \$1779 \$1673 VPWR VGND \$1662 \$1308 VGND
+ sky130_fd_sc_hd__or4_1
X$8610 VPWR \$1783 VPWR VGND \$1649 \$1574 VGND sky130_fd_sc_hd__or2_2
X$8611 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8612 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8613 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8615 VPWR \$1814 VPWR VGND \$1673 \$1532 VGND sky130_fd_sc_hd__or2_2
X$8616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8617 VPWR \$1533 VPWR VGND \$1814 \$1798 VGND sky130_fd_sc_hd__or2_2
X$8618 VPWR \$1801 VPWR VGND \$1574 \$1673 \$1663 VGND sky130_fd_sc_hd__or3_1
X$8619 VPWR VGND VPWR \$1800 \$1706 VGND sky130_fd_sc_hd__inv_2
X$8620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8622 VPWR VGND \$1780 VPWR \$1108 \$1801 VGND sky130_fd_sc_hd__nor2_2
X$8623 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8624 VPWR VGND \$1782 VPWR \$1784 VGND sky130_fd_sc_hd__clkbuf_4
X$8625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8626 VPWR \$1802 \$1707 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8629 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8630 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8631 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8632 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8634 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8635 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8636 VGND \$516 \$1848 \$1273 \$1826 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8638 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8639 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8642 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8643 VGND \$1738 \$1803 mgmt_gpio_out[4] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$8644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8645 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8646 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8647 VPWR \$1760 VGND VPWR \$1767 VGND sky130_fd_sc_hd__clkbuf_1
X$8648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8652 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8654 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8655 VPWR \$2895 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$8656 VPWR VGND irq[1] VPWR \$2895 VGND sky130_fd_sc_hd__buf_2
X$8657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8659 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8660 VPWR \$2997 VGND \$2996 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$8661 VGND \$2997 \$2001 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$8662 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8663 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8664 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8665 VPWR VGND \$2194 VPWR \$2964 VGND sky130_fd_sc_hd__buf_2
X$8666 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8670 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8671 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8672 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8673 VGND \$2930 \$2659 \$2931 \$2942 \$2914 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$8674 VGND \$2659 \$2944 \$2941 \$2893 VPWR \$2990 VPWR VGND
+ sky130_fd_sc_hd__o211ai_4
X$8675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8676 VPWR \$2894 VGND \$2944 VPWR \$2514 VGND sky130_fd_sc_hd__nor2_1
X$8677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8678 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8681 VPWR \$2932 VGND \$2944 VPWR \$2453 VGND sky130_fd_sc_hd__nor2_1
X$8682 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8683 VPWR \$2932 \$2894 VGND \$3054 VPWR \$3011 \$2948 VGND
+ sky130_fd_sc_hd__or4_2
X$8684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8685 VGND \$2946 \$2488 \$2931 \$2943 \$2947 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$8686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8687 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8688 VGND \$2978 \$2949 \$2931 \$2946 \$2965 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$8689 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8691 VPWR VGND VPWR \$2965 \$2797 VGND sky130_fd_sc_hd__inv_2
X$8692 VPWR \$2933 VGND \$2949 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$8693 VPWR \$2797 \$2933 VGND \$2966 VPWR \$2979 \$2948 VGND
+ sky130_fd_sc_hd__or4_2
X$8694 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8696 VPWR VGND VPWR \$2966 \$2951 VGND sky130_fd_sc_hd__inv_2
X$8697 VPWR \$2949 VGND \$2700 \$3958 VPWR \$2952 VGND sky130_fd_sc_hd__o21ai_2
X$8698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8699 VPWR \$2980 VGND \$2933 \$2538 VPWR VGND sky130_fd_sc_hd__or2_1
X$8700 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8701 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8702 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8706 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8707 VGND \$856 \$2859 \$2556 \$2953 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8708 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8709 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8712 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8713 VGND \$856 \$2967 \$2556 \$2981 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8714 VPWR VGND \$2876 \$293 \$2967 \$2981 \$2934 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8716 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8717 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8720 VPWR \$1950 \$2967 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8721 VPWR VGND \$2703 \$281 \$2998 \$3013 \$2705 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8722 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8723 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8724 VGND \$856 \$2935 \$2556 \$2955 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8726 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8727 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8729 VPWR VGND \$1244 VPWR \$2991 \$2897 VGND sky130_fd_sc_hd__nor2_2
X$8730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8731 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8733 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8734 VGND \$2159 \$2956 \$2957 \$2358 \$2274 \$2610 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8735 VGND \$2968 \$2177 \$2983 \$1065 \$880 \$3014 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8736 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8738 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8739 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8740 VGND \$2969 \$1952 \$958 \$2073 \$2096 \$2999 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8741 VPWR VGND VPWR \$2970 \$2969 \$3015 \$2968 \$2042 VGND
+ sky130_fd_sc_hd__and4_1
X$8742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8743 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8744 VGND \$3000 \$3016 \$2593 \$2750 \$2541 \$661 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8746 VPWR \$2984 VGND VPWR \$1097 \$2724 \$2879 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$8747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8749 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8750 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8752 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8753 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8754 VGND \$3001 \$3002 \$2544 \$2545 \$2594 \$2078 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$8755 VGND \$2985 \$2958 \$2594 \$2043 \$1914 \$882 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8757 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8758 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8759 VPWR \$2098 VGND VPWR \$2971 \$2670 \$1817 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$8760 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8761 VPWR \$1490 VGND VPWR \$2325 \$1445 VGND sky130_fd_sc_hd__or2_4
X$8762 VPWR \$1490 VGND VPWR \$2921 \$1426 VGND sky130_fd_sc_hd__or2_4
X$8763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8764 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8765 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8766 VPWR \$1570 VGND VPWR \$2986 \$1454 VGND sky130_fd_sc_hd__or2_4
X$8767 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8768 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8769 VGND \$1105 \$3014 \$2384 \$2162 \$2960 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$8770 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8771 VPWR \$3003 VGND \$1258 \$1571 VPWR VGND sky130_fd_sc_hd__or2_1
X$8772 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8774 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8775 VGND \$3003 \$2919 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$8776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8779 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8781 VGND \$2601 \$3041 \$2807 \$3020 \$2986 \$2992 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$8782 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8783 VPWR \$2987 VGND VPWR \$2917 \$2135 \$2498 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$8784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8785 VGND \$2972 \$2987 \$3004 \$1065 \$880 \$2753 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8786 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8788 VGND \$2961 \$2529 \$2596 \$2073 \$2096 \$2992 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8789 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8791 VPWR VGND VPWR \$2901 \$2961 \$2973 \$2972 \$2588 VGND
+ sky130_fd_sc_hd__and4_1
X$8792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8794 VPWR \$3022 VGND VPWR \$1678 \$1793 \$3005 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$8795 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8797 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8799 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8804 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8806 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8807 VGND \$2865 \$3023 \$500 \$1953 \$1987 \$2403 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8808 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8809 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8810 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8811 VPWR \$2993 VGND VPWR \$1480 \$1793 \$2053 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$8812 VGND \$3025 \$2993 \$2848 \$2065 \$2046 \$2976 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8816 VPWR \$2974 VGND \$2007 \$2880 VPWR VGND sky130_fd_sc_hd__or2_1
X$8817 VGND \$2975 \$2974 \$1521 \$2116 \$1536 \$1221 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$8818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8819 VPWR VGND VPWR \$2905 \$3148 \$2975 \$3056 \$2885 VGND
+ sky130_fd_sc_hd__and4_1
X$8820 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8825 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8826 VGND \$2989 \$2995 \$2450 \$3006 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$8827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8828 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8829 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8830 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8831 VGND \$1152 \$2989 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$8832 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8833 VPWR VGND VPWR \$2694 \$2672 VGND sky130_fd_sc_hd__inv_2
X$8834 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8835 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8837 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8838 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8839 VPWR \$2976 \$2963 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8840 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8841 VPWR VGND \$2730 \$1171 \$3007 \$3027 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$8842 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8844 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8845 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8848 VPWR \$2988 \$2909 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8849 VPWR \$2994 \$3008 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$8850 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8853 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8854 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8856 VPWR VPWR VGND mgmt_gpio_in[8] \$3010 VGND sky130_fd_sc_hd__clkbuf_2
X$8857 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8858 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8861 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8863 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8864 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8865 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8867 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8868 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8870 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8872 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8873 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8874 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8875 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8876 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8878 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8879 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8880 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8882 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8884 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8887 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8888 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8889 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8891 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8892 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8894 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8897 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8898 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8899 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8900 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8901 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8903 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8904 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8905 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8906 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8908 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8910 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8911 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8912 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8913 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8916 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8917 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8918 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8919 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8921 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8923 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8924 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8925 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8926 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8927 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8928 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8930 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8931 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8933 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8934 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8936 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8937 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8938 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8940 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8943 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8944 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8947 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8948 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8949 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8950 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8951 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8952 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8953 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8954 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8955 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8956 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8957 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8959 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8960 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8961 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8962 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8963 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8964 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8965 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8966 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$8968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8969 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8970 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8971 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8972 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8977 VPWR VGND pll_ena VPWR \$194 VGND sky130_fd_sc_hd__buf_2
X$8978 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8979 VGND \$655 \$206 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$8980 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8983 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8984 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$8985 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$8986 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8990 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8992 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8993 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8994 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$8995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8996 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$8997 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$8998 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$8999 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9000 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9001 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9002 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9003 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9004 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9005 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9007 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9008 VPWR \$187 VGND VPWR \$208 VGND sky130_fd_sc_hd__clkbuf_1
X$9009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9011 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9012 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9013 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9014 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9015 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9016 VGND \$206 \$296 \$243 \$209 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9017 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9019 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9020 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9021 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9022 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9023 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9025 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9027 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9028 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9029 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9030 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9031 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9032 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9033 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9035 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9037 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9039 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9040 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9041 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9042 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9043 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9044 VPWR VGND serial_load VPWR \$201 VGND sky130_fd_sc_hd__buf_2
X$9045 VPWR VGND pwr_ctrl_out[2] VPWR \$211 VGND sky130_fd_sc_hd__buf_2
X$9046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9048 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9049 VPWR VGND wb_dat_o[4] VPWR \$4073 VGND sky130_fd_sc_hd__buf_2
X$9050 VPWR VGND wb_dat_o[3] VPWR \$3914 VGND sky130_fd_sc_hd__buf_2
X$9051 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9053 VPWR \$4192 VGND VPWR \$4175 \$3531 \$1975 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$9054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9055 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9056 VPWR \$4137 VGND VPWR \$3470 \$2119 \$2001 \$3833 VGND
+ sky130_fd_sc_hd__o22a_1
X$9057 VGND \$4193 \$3853 \$4176 \$2890 \$4169 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4bb_1
X$9058 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9059 VGND \$4137 \$4169 \$4148 \$3096 VPWR VPWR \$4033 VGND
+ sky130_fd_sc_hd__or4b_1
X$9060 VGND \$4176 \$2537 \$2119 \$4194 \$2336 \$2193 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$9061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9062 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9063 VPWR \$3741 VGND \$4149 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$9064 VPWR \$4177 VGND \$4148 VPWR \$3648 VGND sky130_fd_sc_hd__or2b_1
X$9065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9066 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9067 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9068 VPWR \$4074 VGND \$4113 \$4076 VPWR VGND sky130_fd_sc_hd__or2_1
X$9069 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9071 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9072 VGND \$4048 \$2571 \$3880 \$4177 \$4138 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$9073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9075 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9076 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9077 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9079 VGND \$4178 \$2119 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$9080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9081 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9082 VPWR \$4152 VGND \$4179 VPWR \$4214 VGND sky130_fd_sc_hd__nor2_1
X$9083 VPWR \$4150 VGND \$2472 \$3710 VPWR VGND sky130_fd_sc_hd__or2_1
X$9084 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9085 VPWR \$5350 VPWR VGND \$3700 \$4170 VGND sky130_fd_sc_hd__or2_2
X$9086 VPWR \$4129 \$4150 VPWR \$3710 \$2931 \$4151 VGND \$4139 VGND
+ sky130_fd_sc_hd__o221ai_1
X$9087 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9088 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9089 VPWR \$4196 VPWR VGND \$3652 \$4170 \$4180 VGND sky130_fd_sc_hd__or3b_1
X$9090 VPWR VGND VPWR \$4170 \$4150 VGND sky130_fd_sc_hd__inv_2
X$9091 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9092 VPWR \$4197 VPWR VGND \$4152 \$4140 \$3932 VGND sky130_fd_sc_hd__or3_1
X$9093 VPWR \$4130 VGND \$4129 \$4140 VPWR VGND sky130_fd_sc_hd__or2_1
X$9094 VPWR VGND VPWR \$4114 \$4223 VGND sky130_fd_sc_hd__inv_2
X$9095 VPWR \$4080 VPWR VGND \$4152 \$4114 \$4130 VGND sky130_fd_sc_hd__or3_1
X$9096 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9097 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9098 VPWR \$4153 \$4132 \$4154 VPWR VGND \$4079 \$4131 VGND
+ sky130_fd_sc_hd__or4_1
X$9099 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9100 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9101 VGND \$4156 \$4153 \$4155 \$4141 \$4095 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211ai_2
X$9102 VPWR \$4141 VGND \$4181 VPWR \$4154 VGND sky130_fd_sc_hd__nor2_1
X$9103 VPWR VGND VPWR \$4155 \$4158 VGND sky130_fd_sc_hd__inv_2
X$9104 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9105 VGND \$4157 \$4141 \$4105 \$4133 \$4158 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$9106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9107 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9108 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9112 VPWR VGND VPWR \$3216 \$4198 VGND sky130_fd_sc_hd__inv_2
X$9113 VPWR \$3391 \$4254 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9116 VGND \$2777 \$4171 \$3921 \$4182 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9117 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9118 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9119 VPWR VGND \$4142 VPWR \$4159 \$1341 VGND sky130_fd_sc_hd__nor2_2
X$9120 VPWR VGND VPWR \$4106 \$4142 VGND sky130_fd_sc_hd__inv_4
X$9121 VPWR VGND \$4183 \$4023 \$4184 \$4200 \$4185 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9122 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9123 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9124 VPWR \$4201 VGND \$3181 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$9125 VPWR \$3939 \$4171 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9126 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9128 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9129 VPWR VGND VPWR \$4082 \$4184 VGND sky130_fd_sc_hd__inv_2
X$9130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9131 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9135 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9137 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9138 VGND \$4218 \$4202 \$4023 \$4186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9141 VPWR \$4052 VGND VPWR \$3883 \$2254 \$3939 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$9142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9144 VPWR \$4116 VGND VPWR \$3910 \$2254 \$3999 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$9145 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9146 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9149 VPWR \$4143 VGND VPWR \$3391 \$3703 \$4117 \$3019 VGND
+ sky130_fd_sc_hd__o22a_1
X$9150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9151 VGND \$4160 \$3897 \$3204 \$3019 \$3722 \$3041 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$9152 VPWR \$4160 VGND VPWR \$2900 \$3121 \$3840 \$3703 VGND
+ sky130_fd_sc_hd__o22a_1
X$9153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9155 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9156 VGND \$4025 \$4143 \$3999 \$3181 \$3121 \$4039 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9157 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9158 VGND \$4203 \$4038 \$4082 \$3181 \$2921 \$3979 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9159 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9161 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9162 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9163 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9165 VGND \$4204 \$2249 \$3794 \$2789 \$2031 \$4120 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9167 VPWR \$2249 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9170 VGND \$4256 \$3939 \$3181 \$3765 \$2669 \$2625 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$9171 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9173 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9174 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9175 VGND \$4144 \$4161 \$3768 \$2581 \$2919 \$4110 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9176 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9178 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9179 VPWR \$4121 VGND VPWR \$3746 \$2456 \$4145 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$9180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9182 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9184 VGND \$4205 \$3076 \$2089 \$2073 \$2096 \$4027 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9186 VGND \$4001 \$4206 \$4462 VPWR \$1107 VPWR VGND sky130_fd_sc_hd__nand3_4
X$9187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9189 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9190 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9192 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9195 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9196 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9198 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9199 VGND \$4172 \$4208 \$1077 \$2525 \$2458 \$4187 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9200 VPWR \$1590 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9201 VGND \$3243 \$1590 \$4146 \$2986 \$2614 \$4173 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9203 VGND \$4188 \$4207 \$4030 \$1065 \$880 \$1601 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9205 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9208 VGND \$4162 \$3190 \$4031 \$2073 \$2096 \$4146 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9209 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9210 VPWR VGND VPWR \$4174 \$4162 \$4209 \$4188 \$3687 VGND
+ sky130_fd_sc_hd__and4_1
X$9211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9212 VGND \$4019 \$4174 \$4163 VPWR \$931 VPWR VGND sky130_fd_sc_hd__nand3_4
X$9213 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9214 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9215 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9217 VPWR VGND \$4189 \$2596 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$9218 VGND \$2989 \$4089 \$4164 \$4111 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9220 VGND \$3952 \$4164 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$9221 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9222 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9223 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9224 VPWR VGND \$3717 VPWR \$4135 VGND sky130_fd_sc_hd__clkbuf_4
X$9225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9226 VPWR VGND VPWR \$4085 \$4103 VGND sky130_fd_sc_hd__inv_2
X$9227 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9228 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9230 VPWR VGND \$3716 \$184 \$4091 \$4166 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9231 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9233 VGND \$2989 \$4091 \$4165 \$4166 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9234 VGND \$2989 \$4128 \$4165 \$4136 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$9235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9236 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9237 VGND \$1892 \$4128 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$9238 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9239 VPWR VGND \$3872 \$1594 \$4190 \$4112 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9240 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9241 VGND \$4167 \$2671 mgmt_gpio_out[11] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$9242 VPWR VGND \$4190 \$2669 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$9243 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9244 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9246 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9248 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9251 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9252 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9253 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9254 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9255 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9256 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9257 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9258 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9259 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9260 VPWR \$401 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9261 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9263 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9265 VPWR \$397 VGND VPWR \$359 VGND sky130_fd_sc_hd__clkbuf_1
X$9266 VGND \$376 \$235 \$387 \$408 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$9267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9269 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9270 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9272 VGND \$388 \$308 \$387 \$409 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$9273 VPWR VGND \$428 VPWR \$440 \$308 \$409 VGND sky130_fd_sc_hd__a21o_1
X$9274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9276 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9278 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9279 VPWR \$441 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$9280 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9282 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9283 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9285 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9286 VPWR \$442 \$194 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9287 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9288 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9290 VGND \$206 \$350 \$239 \$444 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9291 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9292 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9293 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9294 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9295 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9296 VGND \$206 \$373 \$239 \$410 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9297 VPWR VGND \$443 \$184 \$373 \$410 \$429 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9299 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9301 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9302 VGND \$206 \$398 \$241 \$423 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9303 VPWR VGND \$204 \$200 \$398 \$423 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9306 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9308 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9309 VPWR VGND \$204 \$411 \$430 \$445 \$205 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9310 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9311 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9314 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9316 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9317 VPWR VGND VPWR \$363 \$346 VGND sky130_fd_sc_hd__inv_2
X$9318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9321 VPWR \$282 \$283 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9322 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9323 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9324 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9326 VPWR VGND \$283 VPWR \$431 VGND sky130_fd_sc_hd__clkbuf_4
X$9327 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9328 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9329 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9331 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9335 VPWR \$413 VGND VPWR \$389 \$325 \$390 \$347 VGND sky130_fd_sc_hd__o22a_1
X$9336 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9337 VGND \$448 \$413 \$424 \$379 \$420 \$364 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9338 VPWR VGND \$230 VPWR \$402 VGND sky130_fd_sc_hd__buf_2
X$9339 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9340 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9341 VPWR \$402 VGND \$420 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$9342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9343 VGND \$432 \$412 \$320 \$433 \$415 \$449 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$9344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9345 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9346 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9347 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9351 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9352 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9354 VGND \$206 \$384 \$243 \$414 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9357 VPWR VGND \$417 \$183 \$384 \$414 \$434 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9359 VPWR VGND VPWR \$390 \$348 VGND sky130_fd_sc_hd__inv_2
X$9360 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9361 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9363 VPWR \$347 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9364 VPWR \$405 VGND \$347 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$9365 VPWR VPWR VGND \$405 \$288 VGND sky130_fd_sc_hd__clkbuf_2
X$9366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9367 VPWR VGND \$271 \$293 \$406 \$416 \$288 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9368 VPWR VGND \$271 \$281 \$399 \$400 \$288 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9369 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9370 VGND \$206 \$406 \$435 \$416 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9372 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9373 VGND \$206 \$399 \$435 \$400 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9375 VPWR VGND VPWR \$417 \$434 VGND sky130_fd_sc_hd__inv_2
X$9376 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9378 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9379 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9380 VGND \$206 \$458 \$435 \$450 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9383 VGND \$422 \$478 \$426 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9384 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9385 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9389 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9390 VGND \$460 \$289 \$436 \$427 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$9391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9393 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9394 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9395 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9398 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9400 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9401 VGND \$418 \$222 \$368 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9403 VGND \$392 \$289 \$393 \$418 \$251 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$9404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9405 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9406 VGND \$206 \$452 \$254 \$419 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9407 VGND \$451 \$452 \$393 \$300 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9408 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9409 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9410 VPWR VGND \$291 \$411 \$452 \$419 \$292 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9411 VGND \$206 \$394 \$254 \$395 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9414 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9415 VGND \$407 \$254 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$9416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9418 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9419 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9420 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9421 VPWR VGND serial_data_2 VPWR \$451 VGND sky130_fd_sc_hd__buf_2
X$9422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9423 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9424 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9426 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9427 VPWR \$718 VGND VPWR sram_ro_data[2] VGND sky130_fd_sc_hd__clkbuf_1
X$9428 VPWR VGND VPWR \$678 \$653 VGND sky130_fd_sc_hd__inv_2
X$9429 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9430 VGND \$679 \$720 \$381 \$719 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$9431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9433 VPWR \$669 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$9434 VPWR \$679 VGND VPWR \$669 VGND sky130_fd_sc_hd__clkbuf_1
X$9435 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9436 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9439 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9442 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9443 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9444 VGND \$680 \$481 \$564 \$597 \$623 \$673 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$9445 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9447 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9448 VPWR VGND VPWR \$673 \$599 VGND sky130_fd_sc_hd__inv_2
X$9449 VPWR \$721 \$700 \$680 \$584 VGND \$709 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$9450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9451 VGND \$813 \$682 \$381 \$700 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9452 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9453 VGND \$600 \$673 \$681 \$682 \$492 VPWR VPWR VGND sky130_fd_sc_hd__a31o_1
X$9454 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9458 VPWR \$722 VGND VPWR \$710 VGND sky130_fd_sc_hd__clkbuf_1
X$9459 VPWR \$710 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$9460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9462 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9463 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9464 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9465 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9466 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9469 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9470 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9473 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9476 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9477 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9478 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9479 VPWR VGND \$701 \$294 \$724 \$723 \$711 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9481 VPWR VGND \$701 \$183 \$641 \$656 \$711 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9482 VPWR VGND VPWR \$701 \$711 VGND sky130_fd_sc_hd__inv_2
X$9483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9484 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9485 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9488 VPWR VGND VPWR \$702 \$641 VGND sky130_fd_sc_hd__inv_2
X$9489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9492 VGND \$655 \$658 \$196 \$657 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9493 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9494 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9495 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9496 VPWR VGND VPWR \$725 \$624 VGND sky130_fd_sc_hd__inv_2
X$9497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9498 VPWR VGND \$514 \$281 \$660 \$659 \$515 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9499 VPWR VGND \$658 \$712 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$9500 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9501 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9502 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9503 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9504 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9505 VGND \$655 \$670 \$196 \$685 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9506 VPWR VGND \$660 \$684 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$9507 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9508 VPWR VGND \$602 \$183 \$670 \$685 \$674 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9510 VPWR VGND VPWR \$602 \$674 VGND sky130_fd_sc_hd__inv_2
X$9511 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9512 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9513 VPWR \$726 \$670 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9514 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9516 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9517 VPWR VPWR VGND \$727 \$568 VGND sky130_fd_sc_hd__clkbuf_2
X$9518 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9519 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9520 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9521 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9522 VPWR VGND \$567 \$293 \$728 \$736 \$568 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9524 VPWR \$703 \$604 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9526 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9528 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9529 VPWR VGND VPWR \$687 \$626 VGND sky130_fd_sc_hd__inv_2
X$9530 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9531 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9533 VGND \$516 \$729 \$605 \$704 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9535 VPWR VGND \$627 \$293 \$729 \$704 \$607 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9537 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9540 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9541 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9542 VPWR VGND VPWR \$688 \$223 VGND sky130_fd_sc_hd__inv_2
X$9543 VGND \$516 \$628 \$435 \$643 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9544 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9545 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9546 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9549 VPWR VGND \$713 \$293 \$730 \$705 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9550 VGND \$516 \$730 \$435 \$705 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9552 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9554 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9555 VGND \$516 \$650 \$435 \$663 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9557 VPWR VGND VPWR \$731 \$650 VGND sky130_fd_sc_hd__inv_2
X$9558 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9559 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9560 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9563 VPWR VGND \$713 \$354 \$690 \$689 \$714 VPWR VGND sky130_fd_sc_hd__a22o_1
X$9564 VGND \$516 \$690 \$435 \$689 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9565 VPWR VGND VPWR \$774 \$690 VGND sky130_fd_sc_hd__inv_2
X$9566 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9567 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9568 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9569 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9570 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9571 VPWR \$675 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9572 VPWR \$675 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9573 VGND \$671 \$690 \$675 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9576 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9577 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9578 VPWR \$691 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9579 VPWR \$691 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9580 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9581 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9582 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9583 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9584 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9585 VGND \$666 \$289 \$665 \$692 \$676 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$9586 VPWR VGND VPWR \$289 \$676 VGND sky130_fd_sc_hd__inv_4
X$9587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9588 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9590 VPWR \$251 VGND VPWR \$715 VGND sky130_fd_sc_hd__buf_1
X$9591 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9592 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9594 VGND \$706 \$289 \$668 \$707 \$716 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$9595 VGND \$206 \$668 \$541 \$706 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9597 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9599 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9600 VGND \$206 \$694 \$541 \$693 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9602 VGND \$693 \$672 \$695 \$677 \$694 \$696 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$9603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9604 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9605 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9606 VGND \$652 \$745 \$698 \$571 \$717 \$677 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$9607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9608 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9609 VGND \$206 \$698 \$541 \$697 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9611 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9612 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9613 VPWR \$732 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9614 VPWR VGND mgmt_gpio_out[0] VPWR \$732 VGND sky130_fd_sc_hd__buf_2
X$9615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9620 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9621 VPWR VGND spi_sdi VPWR \$3388 VGND sky130_fd_sc_hd__buf_2
X$9622 VPWR \$3429 \$3389 VPWR \$3438 VGND VGND sky130_fd_sc_hd__and2_1
X$9623 VPWR \$3388 VGND VPWR \$3389 VGND sky130_fd_sc_hd__clkbuf_1
X$9624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9626 VPWR \$3409 VGND \$2234 VPWR \$3057 VGND sky130_fd_sc_hd__nor2_1
X$9627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9629 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9630 VGND \$3248 \$3341 \$3357 \$3340 \$3409 \$2390 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2111o_1
X$9631 VPWR \$4359 \$3431 \$3430 VPWR VGND \$3357 \$3231 VGND
+ sky130_fd_sc_hd__or4_1
X$9632 VGND \$3341 \$3359 \$3114 \$3410 \$2390 \$3341 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_1
X$9633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9634 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9635 VPWR VGND VPWR \$3359 \$2552 VGND sky130_fd_sc_hd__inv_2
X$9636 VPWR VGND VPWR \$3341 \$3124 VGND sky130_fd_sc_hd__inv_2
X$9637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9639 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9642 VPWR \$2929 \$3432 \$3891 VPWR VGND \$3153 \$3154 VGND
+ sky130_fd_sc_hd__or4_1
X$9643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9645 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9646 VGND \$3453 \$3452 \$3440 \$3439 \$2837 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$9647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9648 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9649 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9651 VPWR \$3441 VGND \$2119 VPWR \$3155 VGND sky130_fd_sc_hd__nor2_1
X$9652 VGND \$3454 \$2156 \$3201 \$3441 \$3442 VPWR VPWR VGND
+ sky130_fd_sc_hd__nor4_2
X$9653 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9654 VPWR \$3412 \$3787 \$2774 VPWR VGND \$3269 \$3453 VGND
+ sky130_fd_sc_hd__or4_1
X$9655 VPWR \$3441 VPWR VGND \$3693 \$3412 \$3433 VGND sky130_fd_sc_hd__or3_2
X$9656 VPWR \$3412 VGND \$3141 VPWR \$1998 VGND sky130_fd_sc_hd__nor2_1
X$9657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9658 VPWR \$3455 VGND \$3178 VPWR \$3412 VGND sky130_fd_sc_hd__nor2_1
X$9659 VPWR \$3433 VGND \$3141 VPWR \$1962 VGND sky130_fd_sc_hd__nor2_1
X$9660 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9663 VPWR \$3456 VGND \$3433 \$3443 VPWR VGND sky130_fd_sc_hd__or2_1
X$9664 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9665 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9666 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9667 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9671 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9672 VPWR VGND VPWR \$3284 \$3304 VGND sky130_fd_sc_hd__inv_2
X$9673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9674 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9675 VGND \$856 \$3414 \$3413 \$3390 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9676 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9677 VPWR VGND \$3284 \$281 \$3414 \$3390 \$3304 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9678 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9680 VGND \$856 \$3345 \$3413 \$3434 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9681 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9682 VPWR \$2593 \$3414 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9683 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9684 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9686 VGND \$856 \$3416 \$3413 \$3415 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9687 VPWR VGND \$3435 \$281 \$3345 \$3434 \$3458 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9688 VPWR VGND \$3435 \$200 \$3416 \$3415 \$3458 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9692 VPWR \$3346 VGND VPWR \$3391 \$2229 \$3307 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$9693 VPWR VGND VPWR \$3307 \$3416 VGND sky130_fd_sc_hd__inv_2
X$9694 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9696 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9697 VPWR \$3347 VGND VPWR \$3392 \$3209 \$1076 \$816 VGND
+ sky130_fd_sc_hd__o22a_1
X$9698 VPWR VGND VPWR \$3392 \$3429 VGND sky130_fd_sc_hd__inv_2
X$9699 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9700 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9701 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9702 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9703 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9704 VPWR \$3445 VGND VPWR \$3444 \$1219 \$815 \$816 VGND
+ sky130_fd_sc_hd__o22a_1
X$9705 VGND \$3393 \$3325 \$3459 VPWR \$619 VPWR VGND sky130_fd_sc_hd__nand3_4
X$9706 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9707 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9708 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9709 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9711 VPWR VGND VPWR \$3393 \$1878 \$3394 \$2061 \$3418 VGND
+ sky130_fd_sc_hd__and4_1
X$9712 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9713 VPWR \$3367 VGND VPWR \$3395 \$1125 \$2609 \$923 VGND
+ sky130_fd_sc_hd__o22a_1
X$9714 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9716 VPWR VGND VPWR \$3419 \$3335 \$3460 \$3203 \$3365 VGND
+ sky130_fd_sc_hd__and4_1
X$9717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9718 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9720 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9722 VGND \$3327 \$3419 \$4040 VPWR \$1829 VPWR VGND sky130_fd_sc_hd__nand3_4
X$9723 VPWR \$572 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9724 VPWR VGND VPWR \$3313 \$3461 \$3366 \$572 \$3370 VGND
+ sky130_fd_sc_hd__and4_1
X$9725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9726 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9727 VPWR \$3369 VGND VPWR \$2804 \$1967 \$2784 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$9728 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9729 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9733 VGND \$3396 \$3328 \$2005 \$3566 \$3371 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$9734 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9735 VGND \$3075 \$3396 \$1025 \$3420 \$3397 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$9736 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9737 VGND \$2727 \$3445 \$3436 \$1125 \$1819 \$3446 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9738 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9739 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9740 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9741 VPWR \$3462 VGND VPWR \$1617 \$1776 \$3364 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$9742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9743 VPWR \$3375 VGND VPWR \$3446 \$2456 \$2992 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$9744 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9745 VGND \$3398 \$3375 \$2917 \$2525 \$2458 \$2853 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9746 VPWR \$3330 VGND VPWR \$3399 \$1967 \$2599 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$9747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9749 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9750 VGND \$3400 \$3463 \$3089 \$2325 \$2447 \$3447 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9751 VPWR \$1509 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9752 VGND \$3421 \$3314 \$1509 \$3400 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$9753 VGND \$3422 \$3378 \$2005 \$3401 \$3377 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$9754 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9755 VGND \$3448 \$3464 \$3422 \$3062 VPWR \$3437 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$9756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9757 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9758 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9759 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9760 VPWR \$1411 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9761 VPWR \$260 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9762 VGND \$3449 \$1411 \$3404 \$2162 \$2497 \$3405 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$9763 VPWR \$3423 VGND VPWR \$3402 \$1645 \$260 \$326 VGND
+ sky130_fd_sc_hd__o22a_1
X$9764 VPWR \$3315 VGND VPWR \$4319 \$1967 \$3403 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$9765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9767 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9768 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9770 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9771 VPWR \$3353 VGND VPWR \$3404 \$1967 \$3405 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$9772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9775 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9776 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9777 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9778 VGND \$3406 \$3424 \$3381 \$3025 VPWR \$675 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$9779 VPWR \$3355 VGND VPWR \$3450 \$2670 \$2630 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$9780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9781 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9782 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9783 VGND \$2989 \$3426 \$3425 \$3407 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9785 VPWR VGND \$2633 \$184 \$3426 \$3407 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9786 VPWR VGND VPWR \$3467 \$3426 VGND sky130_fd_sc_hd__inv_2
X$9787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9788 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9789 VGND \$2989 \$3408 \$3425 \$3427 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9790 VPWR VGND \$2633 \$411 \$3408 \$3427 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9791 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9793 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9794 VPWR VGND \$2694 \$354 \$3428 \$3384 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9795 VPWR VGND VPWR \$3354 \$3428 VGND sky130_fd_sc_hd__inv_2
X$9796 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9797 VPWR \$3378 \$3385 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9798 VGND \$2989 \$3428 \$3425 \$3384 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9799 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9800 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9801 VGND \$2989 \$3385 \$3425 \$3386 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9803 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9804 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9805 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9806 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9808 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9809 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9811 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9812 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9814 VPWR \$3468 VGND VPWR \$2791 VGND sky130_fd_sc_hd__clkbuf_1
X$9815 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9816 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9821 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9822 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9823 VPWR \$1513 \$1522 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9824 VPWR \$1548 \$1577 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9825 VPWR VGND VPWR \$1549 \$1564 VGND sky130_fd_sc_hd__inv_2
X$9826 VPWR \$1522 VGND VPWR sram_ro_data[16] VGND sky130_fd_sc_hd__clkbuf_1
X$9827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9828 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9829 VGND \$1497 \$1186 \$1514 \$1498 \$1523 \$1473 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$9830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9832 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9833 VPWR VGND VPWR \$1514 \$1473 VGND sky130_fd_sc_hd__inv_2
X$9834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9835 VPWR VGND \$1514 \$1524 \$1460 \$1515 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9837 VGND \$864 \$1460 \$387 \$1515 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$9838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9839 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9840 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9841 VPWR \$1565 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$9842 VPWR \$1579 VGND VPWR \$1565 VGND sky130_fd_sc_hd__clkbuf_1
X$9843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9845 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9846 VGND \$1581 \$1433 \$1582 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9847 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9848 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9850 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9851 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9853 VPWR VGND VPWR \$1583 \$1500 VGND sky130_fd_sc_hd__inv_2
X$9854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9855 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9856 VGND \$1687 \$1337 \$1501 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9857 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9858 VGND \$1584 \$1433 \$1580 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9859 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9860 VGND \$1516 \$1487 \$1433 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9861 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9862 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9863 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9865 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9866 VGND \$1474 \$1516 \$1636 \$1369 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$9867 VGND \$1503 \$1550 \$1584 \$1369 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$9868 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9870 VGND \$1503 \$1526 \$1504 \$1525 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$9871 VPWR VGND VPWR \$1504 \$1369 VGND sky130_fd_sc_hd__inv_2
X$9872 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9873 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9874 VGND \$856 \$1540 \$891 \$1539 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9875 VGND \$856 \$1527 \$891 \$1551 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$9876 VPWR VGND \$1399 \$200 \$1527 \$1551 \$1417 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9879 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9880 VPWR VGND \$1399 \$294 \$1566 \$1552 \$1417 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9883 VPWR \$1506 VPWR VGND \$1462 \$1474 \$1526 VGND sky130_fd_sc_hd__or3_1
X$9884 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9885 VPWR \$1517 VPWR VGND \$1462 \$1477 \$1526 VGND sky130_fd_sc_hd__or3_1
X$9886 VPWR \$1553 VPWR VGND \$1477 \$1453 \$1489 VGND sky130_fd_sc_hd__or3_1
X$9887 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9889 VPWR VGND VPWR \$1477 \$1474 VGND sky130_fd_sc_hd__inv_2
X$9890 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9891 VGND \$1517 \$1571 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$9892 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9893 VGND \$1553 \$1570 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$9894 VGND \$856 \$1555 \$922 \$1541 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9895 VPWR \$1542 VGND VPWR \$868 \$1058 \$1549 \$1554 VGND
+ sky130_fd_sc_hd__o22a_1
X$9896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9897 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9898 VPWR VGND \$1567 \$200 \$1555 \$1541 \$1568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9900 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9901 VPWR VGND VPWR \$1569 \$1555 VGND sky130_fd_sc_hd__inv_2
X$9902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9904 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9905 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9906 VPWR \$1444 VGND VPWR \$347 \$1248 VGND sky130_fd_sc_hd__or2_4
X$9907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9908 VPWR \$1435 VGND VPWR \$1554 \$1248 VGND sky130_fd_sc_hd__or2_4
X$9909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9910 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9911 VPWR \$1426 VGND VPWR \$848 \$1248 VGND sky130_fd_sc_hd__or2_4
X$9912 VPWR \$1329 VGND VPWR \$1556 \$1248 VGND sky130_fd_sc_hd__or2_4
X$9913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9915 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9918 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9919 VPWR \$1557 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9920 VPWR \$1585 VGND VPWR \$1350 \$1297 \$1557 \$1219 VGND
+ sky130_fd_sc_hd__o22a_1
X$9921 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9923 VPWR \$1570 VGND VPWR \$1558 \$1434 VGND sky130_fd_sc_hd__or2_4
X$9924 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9925 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9926 VPWR \$1598 VGND VPWR \$859 \$1264 VGND sky130_fd_sc_hd__or2_4
X$9927 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9929 VPWR \$1505 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9930 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9932 VGND \$1508 \$1563 \$848 \$1556 \$1559 \$1560 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$9933 VPWR \$560 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$9934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9935 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9936 VPWR \$1426 VGND VPWR \$1562 \$1571 VGND sky130_fd_sc_hd__or2_4
X$9937 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9938 VPWR \$1445 VGND VPWR \$1465 \$1248 VGND sky130_fd_sc_hd__or2_4
X$9939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9940 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9941 VPWR \$1454 VGND VPWR \$1561 \$1571 VGND sky130_fd_sc_hd__or2_4
X$9942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9943 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9944 VPWR \$1528 VGND \$1558 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$9945 VPWR VPWR VGND \$1528 \$1166 VGND sky130_fd_sc_hd__clkbuf_2
X$9946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9947 VPWR VGND VPWR \$1968 \$1455 VGND sky130_fd_sc_hd__inv_2
X$9948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9950 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9951 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9952 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9953 VPWR \$1529 \$1467 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$9954 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9955 VGND \$1152 \$1591 \$771 \$1573 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$9959 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9963 VPWR VGND \$1303 \$200 \$1518 \$1456 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9965 VPWR VGND VPWR \$1617 \$1518 VGND sky130_fd_sc_hd__inv_2
X$9966 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9968 VGND \$1152 \$1530 \$1203 \$1543 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9969 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9971 VPWR VGND \$1303 \$411 \$1530 \$1543 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9973 VPWR VPWR VGND \$1446 \$358 VGND sky130_fd_sc_hd__clkbuf_2
X$9974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9976 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9977 VPWR VGND \$1170 \$200 \$1604 \$1586 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9978 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$9981 VPWR VGND \$1170 \$354 \$1519 \$1544 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$9982 VGND \$1152 \$1519 \$1203 \$1544 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$9983 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$9984 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9986 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9989 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9990 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$9991 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$9993 VPWR \$1011 \$1510 \$1531 \$1545 VGND \$1532 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$9994 VPWR VGND VPWR \$1532 \$1574 VGND sky130_fd_sc_hd__inv_2
X$9995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$9996 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9997 VPWR VGND \$1533 VPWR \$895 \$1545 \$672 VGND sky130_fd_sc_hd__a21oi_1
X$9998 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$9999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10000 VGND \$1520 \$1534 \$1470 \$1535 \$1536 \$1011 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$10001 VPWR \$1533 \$1535 VGND \$1011 VPWR \$1575 VGND sky130_fd_sc_hd__nor3_1
X$10002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10003 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10004 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10005 VPWR \$1537 \$1535 VPWR \$1545 VGND \$1546 VGND sky130_fd_sc_hd__o21ba_1
X$10006 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10007 VGND \$516 \$1546 \$541 \$1537 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10008 VPWR VGND VPWR \$1534 \$1576 VGND sky130_fd_sc_hd__inv_2
X$10009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10011 VGND \$516 \$1482 \$1273 \$1511 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10013 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10014 VGND \$732 \$1482 \$839 \$1587 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$10015 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10016 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10017 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10018 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10019 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10021 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10022 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10023 VGND \$1512 \$1521 mgmt_gpio_out[3] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$10024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10025 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10026 VPWR \$1471 VGND VPWR \$1521 VGND sky130_fd_sc_hd__clkbuf_1
X$10027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10030 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10031 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10032 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10033 VGND \$4862 \$4651 \$5153 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$10034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10037 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10039 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10041 VPWR \$5025 \$5154 \$4942 VPWR VGND \$4941 \$5147 VGND
+ sky130_fd_sc_hd__or4_1
X$10042 VPWR \$4930 \$5155 \$4942 VPWR VGND \$4941 \$5147 VGND
+ sky130_fd_sc_hd__or4_1
X$10043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10044 VGND \$5155 \$2996 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$10045 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10046 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10048 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10049 VGND \$5124 \$5169 \$4891 \$4880 \$4853 \$5181 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$10050 VPWR \$4891 VGND \$5169 \$5089 VPWR \$5181 VGND sky130_fd_sc_hd__o21ai_2
X$10051 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10052 VPWR \$5139 VPWR VGND \$5169 \$5170 \$4854 VGND sky130_fd_sc_hd__or3b_1
X$10053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10055 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10057 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10058 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10061 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10062 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10063 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10064 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10065 VGND \$1897 \$4153 \$4673 VPWR VPWR VGND sky130_fd_sc_hd__nor2_4
X$10066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10067 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10068 VPWR \$5183 VGND \$4737 \$4736 VPWR VGND sky130_fd_sc_hd__or2_1
X$10069 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10070 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10071 VPWR \$5174 VGND \$5233 \$4737 VPWR VGND sky130_fd_sc_hd__or2_1
X$10072 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10073 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10076 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10077 VPWR \$5171 VPWR VGND \$4676 \$4727 \$5174 VGND sky130_fd_sc_hd__or3_1
X$10078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10079 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10080 VPWR \$5247 VGND \$4954 \$4665 VPWR VGND sky130_fd_sc_hd__or2_1
X$10081 VPWR \$5175 VGND \$5171 VPWR \$4954 VGND sky130_fd_sc_hd__nor2_1
X$10082 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10084 VPWR \$5029 VGND \$5246 \$5175 VPWR VGND sky130_fd_sc_hd__or2_1
X$10085 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10086 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10087 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10088 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10090 VPWR \$5163 VGND \$5184 VPWR \$5149 VGND sky130_fd_sc_hd__nor2_1
X$10091 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10092 VPWR VGND VPWR \$5184 \$1315 VGND sky130_fd_sc_hd__inv_2
X$10093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10096 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10097 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10099 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10101 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10102 VGND \$4761 \$5156 \$5165 \$5164 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10103 VPWR VGND \$5118 \$3732 \$5156 \$5164 \$5080 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10104 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10105 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10107 VGND \$4761 \$5158 \$5165 \$5157 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10108 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10113 VGND \$4761 \$5166 \$4813 \$5172 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10115 VPWR \$4117 \$5166 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10117 VPWR VGND \$5086 \$3711 \$5166 \$5172 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10118 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10120 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10122 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10123 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10125 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10126 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10127 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10131 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10133 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10135 VGND \$4761 \$5150 \$4850 \$5142 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10136 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10137 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10138 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10140 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10141 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10146 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10147 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10150 VGND \$4764 \$5151 \$5006 \$5159 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10151 VPWR VGND \$5086 \$411 \$5151 \$5159 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10153 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10154 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10157 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10161 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10162 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10163 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10164 VGND \$4764 \$5160 \$5006 \$5143 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10167 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10169 VPWR \$3092 \$5160 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$10170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10174 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10175 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10176 VPWR VGND \$5046 \$3694 \$5177 \$5173 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10180 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10181 VPWR \$2880 \$5177 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$10182 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10183 VPWR user_clock VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10185 VGND \$5136 user_clock \$5122 \$5068 VPWR VPWR VGND
+ sky130_fd_sc_hd__mux2_1
X$10186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10188 VPWR VGND \$4650 \$354 \$5161 \$5188 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10190 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10192 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10193 VGND \$4764 \$5162 \$4828 \$5168 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10194 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10195 VPWR VGND \$4650 \$1594 \$5162 \$5168 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10196 VPWR VGND VPWR \$4650 \$4659 VGND sky130_fd_sc_hd__inv_2
X$10197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10198 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10199 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10201 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10202 VPWR VGND VPWR \$4236 \$5178 VGND sky130_fd_sc_hd__inv_2
X$10203 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10204 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10205 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10209 VPWR VGND irq[2] VPWR \$2991 VGND sky130_fd_sc_hd__buf_2
X$10210 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10212 VPWR \$2991 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10213 VGND \$1979 \$3067 \$3057 \$2015 VPWR VPWR VGND sky130_fd_sc_hd__nor3_2
X$10214 VPWR \$2015 \$3068 VGND \$3057 VPWR \$1962 VGND sky130_fd_sc_hd__nor3_1
X$10215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10218 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10220 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10222 VPWR \$3069 VGND \$2891 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$10223 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10225 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10226 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10228 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10229 VPWR \$3054 \$3058 VPWR \$2659 \$2944 \$2944 VGND \$2891 VGND
+ sky130_fd_sc_hd__o221ai_1
X$10230 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10231 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10233 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10234 VPWR VGND \$2453 VPWR \$3029 VGND sky130_fd_sc_hd__buf_2
X$10235 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10236 VPWR VGND VPWR \$2224 \$2996 VGND sky130_fd_sc_hd__inv_2
X$10237 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10241 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10246 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10247 VPWR VGND VPWR \$2775 \$2776 VGND sky130_fd_sc_hd__inv_2
X$10248 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10249 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10250 VGND \$2777 \$3012 \$2556 \$3055 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10251 VPWR VGND \$2775 \$281 \$3012 \$3055 \$2776 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10252 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10253 VPWR VPWR VGND \$3059 \$2776 VGND sky130_fd_sc_hd__clkbuf_2
X$10254 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10255 VPWR \$2879 \$3012 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10257 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10258 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10259 VGND \$3030 \$2556 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$10260 VPWR \$3059 VGND \$2372 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$10261 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10264 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10265 VGND \$856 \$2998 \$2556 \$3013 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10268 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10269 VPWR VGND VPWR \$3014 \$2998 VGND sky130_fd_sc_hd__inv_2
X$10270 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10272 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10274 VGND \$3015 \$3031 \$2382 \$2330 \$2219 \$2982 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10276 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10279 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10280 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10282 VPWR \$3016 VGND VPWR \$958 \$2559 \$3017 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$10283 VGND \$3032 \$2984 \$684 \$2369 \$2357 \$2983 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10284 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10285 VGND \$3018 \$2970 \$3033 VPWR \$540 VPWR VGND sky130_fd_sc_hd__nand3_4
X$10286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10287 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10288 VGND \$3000 \$3073 \$2064 \$3032 \$3072 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$10289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10290 VPWR VGND VPWR \$3018 \$1938 \$3034 \$2985 \$3040 VGND
+ sky130_fd_sc_hd__and4_1
X$10291 VPWR \$3001 VGND VPWR \$3035 \$2665 \$3014 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$10292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10294 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10295 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10296 VPWR \$1570 VGND VPWR \$3019 \$1445 VGND sky130_fd_sc_hd__or2_4
X$10297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10299 VPWR \$1235 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10300 VPWR \$3074 VGND VPWR \$1383 \$1776 \$1235 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$10301 VPWR \$4000 VGND VPWR \$1529 \$1558 \$2988 \$2785 VGND
+ sky130_fd_sc_hd__o22a_1
X$10302 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10303 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10304 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10305 VPWR \$3060 VGND \$1445 \$1571 VPWR VGND sky130_fd_sc_hd__or2_1
X$10306 VGND \$3060 \$4239 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$10307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10309 VPWR \$3043 VGND VPWR \$1383 \$1793 \$2191 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$10310 VGND \$3075 \$3043 \$2464 \$2065 \$2046 \$3061 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10312 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10313 VPWR \$3020 VGND VPWR \$2748 \$3106 \$3004 \$2918 VGND
+ sky130_fd_sc_hd__o22a_1
X$10314 VPWR VGND VPWR \$3087 \$3077 \$3046 \$3088 \$2959 VGND
+ sky130_fd_sc_hd__and4_1
X$10315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10318 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10319 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10320 VPWR \$3076 VGND VPWR \$758 \$2045 \$2988 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$10321 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10322 VPWR \$3021 VGND VPWR \$1617 \$1793 \$1915 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$10323 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10324 VGND \$3044 \$3021 \$2449 \$2065 \$2046 \$2988 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10325 VGND \$3062 \$3022 \$2252 \$2065 \$2046 \$2994 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10326 VPWR \$3045 VGND VPWR \$1225 \$2180 \$2982 \$3042 VGND
+ sky130_fd_sc_hd__o22a_1
X$10327 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10328 VPWR \$2474 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10330 VGND \$3046 \$2962 \$3036 \$3019 \$2581 \$2791 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10331 VGND \$3077 \$3045 \$3063 \$2474 \$2921 \$2829 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10332 VPWR \$3078 VGND VPWR \$2432 \$1956 \$1802 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$10333 VPWR \$3047 VGND VPWR \$1603 \$1793 \$1802 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$10334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10335 VGND \$3064 \$3047 \$1823 \$2065 \$2046 \$2813 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10336 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10337 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10339 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10340 VPWR \$3023 VGND VPWR \$2960 \$1967 \$3037 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$10341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10344 VPWR \$3024 VGND VPWR \$1720 \$1793 \$2307 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$10345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10346 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10347 VGND \$3048 \$3024 \$2548 \$2065 \$2046 \$3038 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10351 VGND \$3056 \$3065 \$2908 \$2043 \$1914 \$1803 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10354 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10357 VGND \$1152 \$3049 \$2450 \$3039 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10358 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10359 VPWR VGND \$2401 \$184 \$3049 \$3039 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10361 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10362 VPWR \$3089 \$2995 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10365 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10366 VPWR VGND \$2401 \$386 \$2995 \$3006 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10367 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10369 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10371 VGND \$2989 \$3050 \$2450 \$3026 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10372 VPWR VGND \$2694 \$184 \$3050 \$3026 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10374 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10375 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10377 VPWR VGND VPWR \$3061 \$3007 VGND sky130_fd_sc_hd__inv_2
X$10378 VGND \$2989 \$3007 \$2450 \$3027 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10380 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10381 VPWR VGND VPWR \$3038 \$3051 VGND sky130_fd_sc_hd__inv_2
X$10382 VGND \$2989 \$3051 \$2232 \$3052 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10383 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10384 VPWR VGND \$2730 \$184 \$3051 \$3052 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10385 VPWR VGND \$2730 \$1179 \$3008 \$3053 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10386 VGND \$1152 \$3008 \$2232 \$3053 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10388 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10389 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10391 VPWR \$3079 VGND VPWR \$3066 VGND sky130_fd_sc_hd__clkbuf_1
X$10392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10393 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10398 VPWR uart_enabled VPWR VGND \$2551 VGND sky130_fd_sc_hd__buf_4
X$10399 VGND spi_enabled \$3438 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$10400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10402 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10404 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10405 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10406 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10407 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10408 VPWR \$3661 \$3594 \$3699 VPWR VGND \$3649 \$3616 VGND
+ sky130_fd_sc_hd__or4_1
X$10409 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10410 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10411 VGND \$3690 \$3662 \$3125 \$3680 \$3689 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4bb_1
X$10412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10413 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10414 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10416 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10417 VPWR \$3690 VGND \$3124 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$10418 VGND \$3638 \$3651 \$3691 \$3690 \$3742 \$2571 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$10419 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10420 VPWR \$3651 VGND \$2931 \$3124 VPWR VGND sky130_fd_sc_hd__or2_1
X$10421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10423 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10424 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10426 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10427 VPWR \$3692 VGND \$1897 \$3709 VPWR VGND sky130_fd_sc_hd__or2_1
X$10428 VGND \$3692 \$3639 \$3442 \$3693 VPWR VPWR \$3700 VGND
+ sky130_fd_sc_hd__or4b_1
X$10429 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10430 VPWR \$3701 VPWR VGND \$3692 \$3504 VGND sky130_fd_sc_hd__nand2_1
X$10431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10432 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10433 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10434 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10435 VPWR \$3474 VGND \$3710 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$10436 VPWR \$3572 VGND \$2511 VPWR \$3710 VGND sky130_fd_sc_hd__nor2_1
X$10437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10439 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10441 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10442 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10443 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10444 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10445 VGND \$2777 \$3668 \$3413 \$3683 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10447 VPWR VGND \$3667 \$293 \$3684 \$3731 \$3669 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10448 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10449 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10451 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10452 VGND \$2777 \$2877 \$3413 \$3685 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10455 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10456 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10458 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10459 VGND \$3711 \$200 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$10460 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10461 VPWR VPWR VGND \$3363 \$3702 VGND sky130_fd_sc_hd__clkbuf_2
X$10462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10465 VGND \$3694 \$281 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$10466 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10468 VPWR \$1570 VGND VPWR \$3703 \$1257 VGND sky130_fd_sc_hd__or2_4
X$10469 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10470 VPWR \$2279 VGND VPWR \$3712 \$2229 \$3719 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$10471 VPWR \$1257 VGND VPWR \$3209 \$1571 VGND sky130_fd_sc_hd__or2_4
X$10472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10473 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10476 VGND \$2645 \$2896 \$3553 \$3143 \$3713 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$10477 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10479 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10480 VPWR \$3695 VGND VPWR \$3564 \$2927 \$1115 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$10481 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10483 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10484 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10485 VGND \$2479 \$3695 \$3704 \$2830 \$2651 \$3643 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10488 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10490 VPWR \$3720 VGND VPWR \$1080 \$1558 \$3704 \$3204 VGND
+ sky130_fd_sc_hd__o22a_1
X$10491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10492 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10495 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10497 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10498 VPWR \$3705 VGND VPWR \$1678 \$1776 \$3312 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$10499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10500 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10504 VGND \$3706 \$3705 \$2790 \$1715 \$1754 \$1030 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10506 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10507 VPWR \$3724 VGND VPWR \$3722 \$2229 \$3436 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$10508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10511 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10512 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10513 VGND \$2973 \$3724 \$3723 \$2330 \$2219 \$2647 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10514 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10517 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10518 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10519 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10520 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10522 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10524 VPWR \$3726 VGND VPWR \$1603 \$1776 \$3714 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$10525 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10526 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10527 VGND \$3707 \$3715 \$1603 \$1300 \$1219 \$3714 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10531 VPWR \$1428 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10532 VPWR VGND VPWR \$3728 \$1428 \$2482 \$3727 \$3707 VGND
+ sky130_fd_sc_hd__and4_1
X$10533 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10535 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10536 VPWR \$3708 VGND VPWR \$1390 \$2724 \$2628 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$10537 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10540 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10542 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10545 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10546 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10548 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10549 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10550 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10554 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10555 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10558 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10559 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10560 VPWR VGND \$3716 \$354 \$3730 \$3729 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10561 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10563 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10565 VPWR VGND VPWR \$2806 \$3697 VGND sky130_fd_sc_hd__inv_2
X$10566 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10567 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10568 VGND \$2989 \$3697 \$3590 \$3718 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10569 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10570 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10572 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10575 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10576 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10577 VGND \$3870 mgmt_gpio_in[10] VPWR VPWR VGND
+ sky130_fd_sc_hd__dlymetal6s2s_1
X$10578 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10580 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10584 VPWR VGND irq[0] VPWR \$2733 VGND sky130_fd_sc_hd__buf_2
X$10585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10587 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10588 VPWR VGND \$2537 VPWR \$2890 \$2234 VGND sky130_fd_sc_hd__nor2_2
X$10589 VPWR \$2911 VGND \$2833 \$2890 VPWR VGND sky130_fd_sc_hd__or2_1
X$10590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10592 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10593 VPWR \$2870 VGND \$2472 VPWR \$2891 VGND sky130_fd_sc_hd__nor2_1
X$10594 VPWR \$2939 VGND \$2890 \$2912 VPWR VGND sky130_fd_sc_hd__or2_1
X$10595 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10596 VPWR \$2892 \$2658 \$2912 VPWR VGND \$2870 \$2835 VGND
+ sky130_fd_sc_hd__or4_1
X$10597 VPWR \$2912 VGND \$2511 VPWR \$2891 VGND sky130_fd_sc_hd__nor2_1
X$10598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10599 VPWR \$2835 VGND \$2891 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$10600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10601 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10602 VPWR VGND \$2925 \$2913 \$2929 VPWR \$2940 \$2195 VGND
+ sky130_fd_sc_hd__or4b_2
X$10603 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10604 VPWR VGND VPWR \$2913 \$2858 VGND sky130_fd_sc_hd__inv_2
X$10605 VPWR \$2914 VGND \$2835 VPWR \$2913 VGND sky130_fd_sc_hd__nor2_1
X$10606 VPWR \$2741 \$2925 \$2891 \$2001 VGND \$2194 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$10607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10608 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10609 VGND \$2941 \$2914 \$2698 \$2816 \$2944 \$2891 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$10610 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10611 VPWR \$2872 VGND \$2521 VPWR \$2795 VGND sky130_fd_sc_hd__nor2_1
X$10612 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10613 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10614 VGND \$2893 \$2552 \$2514 \$2661 \$2872 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$10615 VGND \$2926 \$2514 \$2931 \$2930 \$2872 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$10616 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10617 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10618 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10619 VPWR VGND VPWR \$2915 \$2715 VGND sky130_fd_sc_hd__inv_2
X$10620 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10621 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10622 VPWR \$2715 \$2391 VGND \$2836 VPWR \$2873 \$2894 VGND
+ sky130_fd_sc_hd__or4_2
X$10623 VGND \$2943 \$2453 \$2931 \$2926 \$2915 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$10624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10625 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10626 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10627 VPWR \$2932 \$2796 VGND \$2642 VPWR \$2945 \$2873 VGND
+ sky130_fd_sc_hd__or4_2
X$10628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10629 VPWR VGND VPWR \$2947 \$2642 VGND sky130_fd_sc_hd__inv_2
X$10630 VPWR \$2948 VGND \$2944 VPWR \$2488 VGND sky130_fd_sc_hd__nor2_1
X$10631 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10633 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10634 VPWR \$2950 VGND \$2173 \$2933 VPWR VGND sky130_fd_sc_hd__or2_1
X$10635 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10636 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10637 VPWR \$2774 VGND \$2949 VPWR \$2742 VGND sky130_fd_sc_hd__nor2_1
X$10638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10639 VPWR \$2951 VGND \$2949 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$10640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10641 VPWR \$2798 \$2952 VPWR \$2951 VGND VGND sky130_fd_sc_hd__and2_1
X$10642 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10643 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10644 VGND \$2777 \$2875 \$2556 \$2851 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10647 VPWR \$2383 \$2875 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10648 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10649 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10650 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10652 VPWR VGND \$2876 \$183 \$2859 \$2953 \$2934 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10654 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10655 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10656 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10657 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10658 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10661 VPWR VPWR VGND \$2954 \$1902 VGND sky130_fd_sc_hd__clkbuf_2
X$10662 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10664 VPWR VGND \$2703 \$294 \$2935 \$2955 \$2705 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10665 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10667 VPWR VGND VPWR \$2916 \$2455 VGND sky130_fd_sc_hd__inv_2
X$10668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10669 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10670 VPWR VGND \$1232 VPWR \$2895 \$2756 VGND sky130_fd_sc_hd__nor2_2
X$10671 VPWR VGND VPWR \$2781 \$2935 VGND sky130_fd_sc_hd__inv_2
X$10672 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10674 VPWR \$2956 VGND VPWR \$2383 \$1954 \$2936 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$10675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10677 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10678 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10681 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10682 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10683 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10684 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10685 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10686 VPWR \$2861 VGND VPWR \$2896 \$2665 \$2781 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$10687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10688 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10689 VPWR \$2958 VGND VPWR \$2916 \$1966 \$1948 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$10690 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10691 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10692 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10693 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10694 VPWR \$2562 VGND VPWR \$2917 \$1089 \$2780 \$2314 VGND
+ sky130_fd_sc_hd__o22a_1
X$10695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10696 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10697 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10698 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10699 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10700 VPWR \$1570 VGND VPWR \$2918 \$1329 VGND sky130_fd_sc_hd__or2_4
X$10701 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10702 VPWR \$1490 VGND VPWR \$2180 \$1454 VGND sky130_fd_sc_hd__or2_4
X$10703 VPWR \$1891 VGND VPWR \$2879 \$2372 \$2854 \$2375 VGND
+ sky130_fd_sc_hd__o22a_1
X$10704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10705 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10706 VPWR \$2920 VGND VPWR \$2898 \$2919 \$661 \$1507 VGND
+ sky130_fd_sc_hd__o22a_1
X$10707 VGND \$2959 \$2920 \$2916 \$2190 \$2918 \$2862 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10709 VPWR VGND VPWR \$2898 \$1424 VGND sky130_fd_sc_hd__inv_2
X$10710 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10711 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10712 VPWR \$1060 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10713 VPWR \$2899 VGND VPWR \$762 \$1060 \$2853 \$2921 VGND
+ sky130_fd_sc_hd__o22a_1
X$10714 VGND \$2565 \$2899 \$2603 \$1879 \$2919 \$2897 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10717 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10718 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10719 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10720 VGND \$2844 \$2901 \$2902 VPWR \$1063 VPWR VGND sky130_fd_sc_hd__nand3_4
X$10721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10723 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10724 VPWR \$1060 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$10725 VPWR \$2962 VGND VPWR \$2923 \$2031 \$882 \$1060 VGND
+ sky130_fd_sc_hd__o22a_1
X$10726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10727 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10729 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10731 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10732 VPWR \$2922 VGND VPWR \$3036 \$2927 \$1925 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$10733 VGND \$2811 \$2922 \$2880 \$2830 \$2651 \$2906 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10735 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10736 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10738 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10739 VPWR \$2928 VGND VPWR \$1373 \$2135 \$2960 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$10740 VGND \$2883 \$2928 \$2862 \$1065 \$880 \$2111 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10745 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10748 VPWR VGND VPWR \$2904 \$2884 \$2903 \$2883 \$2812 VGND
+ sky130_fd_sc_hd__and4_1
X$10749 VGND \$2905 \$2904 \$2907 VPWR \$1036 VPWR VGND sky130_fd_sc_hd__nand3_4
X$10750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10751 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10752 VPWR \$2867 VGND VPWR \$2906 \$2254 \$2866 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$10753 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10754 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10755 VPWR VGND VPWR \$2841 \$2868 VGND sky130_fd_sc_hd__inv_2
X$10756 VGND \$1152 \$2868 \$2450 \$2886 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10757 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10758 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10759 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10760 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10761 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10763 VGND \$2908 \$2855 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$10764 VGND \$2937 \$2450 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$10765 VGND \$1152 \$2832 \$2450 \$2888 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10766 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10768 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10770 VPWR VGND \$2730 \$354 \$2963 \$2889 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10773 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10776 VGND \$1152 \$2909 \$2232 \$2938 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10777 VPWR VGND \$2730 \$386 \$2909 \$2938 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10778 VGND \$1895 \$2906 mgmt_gpio_out[7] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$10779 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10781 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10782 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10783 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10784 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10786 VGND \$1207 \$945 \$381 \$1185 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10787 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10788 VPWR \$1207 VGND VPWR \$1213 VGND sky130_fd_sc_hd__clkbuf_1
X$10789 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10790 VPWR \$1213 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$10791 VPWR \$1185 VGND VPWR \$1143 VGND sky130_fd_sc_hd__clkbuf_1
X$10792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10794 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10795 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10796 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10797 VGND \$1102 \$790 \$828 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$10798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10799 VGND \$1187 \$1188 \$623 \$1069 \$801 \$790 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$10800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10801 VPWR VGND \$733 \$1186 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$10802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10804 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10806 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10807 VPWR \$1214 VGND \$623 VPWR \$564 VGND sky130_fd_sc_hd__nor2_1
X$10808 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10809 VPWR \$1227 VGND VPWR \$428 \$1214 \$1215 \$1208 VGND
+ sky130_fd_sc_hd__o22a_1
X$10810 VPWR \$1208 VGND \$428 VPWR \$1042 VGND sky130_fd_sc_hd__nor2_1
X$10811 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10812 VPWR \$1228 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$10813 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10814 VGND \$1245 \$1162 \$387 \$1189 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$10815 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10816 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10817 VPWR VGND \$1053 \$1174 \$1162 \$1189 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10819 VPWR \$1190 \$1162 VPWR \$1162 VGND \$1145 \$1145 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$10820 VGND \$1174 \$1002 \$1190 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$10821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10822 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10823 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10824 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10825 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10826 VGND \$1229 \$1002 \$1162 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$10827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10828 VGND \$1191 \$986 \$1002 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$10829 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10830 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10831 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10832 VGND \$856 \$1146 \$891 \$1147 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10833 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10834 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10835 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10836 VGND \$463 \$891 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$10837 VPWR VGND \$1087 \$281 \$1231 \$1209 \$1088 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10838 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10839 VPWR VGND \$1087 \$294 \$1216 \$1210 \$1088 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10841 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10842 VGND \$856 \$1216 \$891 \$1210 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10844 VPWR VGND VPWR \$1192 \$1094 VGND sky130_fd_sc_hd__inv_2
X$10845 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10847 VGND \$856 \$1233 \$922 \$1193 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10848 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10850 VPWR \$1193 VGND VPWR \$1175 VGND sky130_fd_sc_hd__clkbuf_1
X$10851 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10852 VGND \$856 \$1194 \$922 \$1148 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10853 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10854 VGND \$1133 \$1194 \$293 \$1217 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$10855 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10857 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10858 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10859 VPWR \$1217 VGND \$1218 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$10860 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10861 VPWR \$1244 \$1194 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10862 VGND \$655 \$1195 \$961 \$1165 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10863 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10864 VGND \$1234 \$1244 \$1218 \$320 \$315 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$10865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10866 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10868 VPWR VGND \$892 \$200 \$1195 \$1165 \$911 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10869 VGND \$655 \$1176 \$961 \$1196 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10870 VPWR VGND \$892 \$183 \$1176 \$1196 \$911 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10871 VPWR VPWR VGND \$1149 \$911 VGND sky130_fd_sc_hd__clkbuf_2
X$10872 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10873 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10874 VPWR \$1236 \$1176 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10875 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10876 VPWR \$1197 VGND VPWR \$442 \$353 \$1071 \$1198 VGND
+ sky130_fd_sc_hd__o22a_1
X$10877 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10878 VGND \$1220 \$1197 \$1235 \$1219 \$566 \$1164 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10880 VGND \$1199 \$1150 \$702 \$1058 \$755 \$267 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10882 VPWR VGND VPWR \$1238 \$1199 \$1220 \$1237 \$448 VGND
+ sky130_fd_sc_hd__and4_1
X$10883 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10884 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10885 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10886 VGND \$655 \$1177 \$605 \$1200 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10887 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10888 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10889 VPWR VGND \$912 \$183 \$1177 \$1200 \$893 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10890 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10894 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10896 VPWR \$319 VPWR VGND \$1420 \$1248 VGND sky130_fd_sc_hd__or2_2
X$10897 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10898 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10899 VPWR VGND \$1178 \$1179 \$1151 \$1126 \$1166 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10900 VPWR VGND VPWR \$1239 \$1151 VGND sky130_fd_sc_hd__inv_2
X$10901 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10902 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10903 VPWR VGND \$1178 \$294 \$1167 \$1168 \$1166 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10904 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10905 VPWR \$1240 \$1167 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10906 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10908 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10909 VGND \$1152 \$1167 \$771 \$1168 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10911 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10912 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10913 VPWR \$1202 \$1153 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$10914 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10915 VGND \$655 \$1153 \$1203 \$1154 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10920 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10921 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10922 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10923 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10924 VGND \$1180 \$1047 \$1169 \$1156 \$1157 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$10925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10926 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10927 VPWR VGND VPWR \$1181 \$1071 VGND sky130_fd_sc_hd__inv_4
X$10928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10929 VPWR VGND \$1170 \$1171 \$1181 \$1204 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10930 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10931 VGND \$516 \$1181 \$993 \$1204 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$10932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10933 VPWR VGND \$1170 \$281 \$1172 \$1158 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$10934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$10935 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10936 VGND \$1221 \$1172 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$10937 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10938 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10940 VGND \$516 \$1138 \$1201 \$1173 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10941 VPWR \$1159 VPWR \$1173 VGND \$1205 \$1222 VGND sky130_fd_sc_hd__o21a_1
X$10942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10943 VGND \$1211 \$895 \$1212 \$1260 \$1223 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$10944 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10945 VGND \$516 \$1137 \$1201 \$1211 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$10946 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10947 VGND \$1223 \$1011 \$1128 \$1205 \$1137 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$10948 VPWR VGND VPWR \$1212 \$1128 VGND sky130_fd_sc_hd__inv_2
X$10949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10950 VGND \$1160 \$1183 \$1171 \$520 \$560 \$1129 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10952 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10953 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10954 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10955 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10956 VGND \$516 \$1139 \$466 \$1161 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$10957 VPWR \$1205 VPWR VGND \$895 \$1184 VGND sky130_fd_sc_hd__or2_2
X$10958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10959 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$10960 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10961 VGND \$1141 \$1139 \$914 \$1012 \$1184 \$745 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$10962 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10963 VGND \$1309 \$1140 \$914 \$1012 \$1142 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2bb2o_1
X$10964 VPWR VGND VPWR \$1184 \$1140 VGND sky130_fd_sc_hd__inv_2
X$10965 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10966 VPWR VGND VPWR \$1142 \$1129 VGND sky130_fd_sc_hd__inv_2
X$10967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10968 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10969 VGND \$358 \$407 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$10970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10971 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10975 VGND mgmt_gpio_in[2] \$780 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$10976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10977 VPWR \$1241 VGND VPWR \$1224 VGND sky130_fd_sc_hd__clkbuf_1
X$10978 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10979 VPWR \$1224 VGND VPWR \$1225 VGND sky130_fd_sc_hd__clkbuf_1
X$10980 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10981 VPWR VGND mgmt_gpio_oeb[2] VPWR \$1241 VGND sky130_fd_sc_hd__buf_2
X$10982 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10983 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10984 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10985 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$10986 VPWR VGND wb_dat_o[15] VPWR \$4696 VGND sky130_fd_sc_hd__buf_2
X$10987 VGND \$4438 \$4651 \$4732 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$10988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10989 VPWR \$4732 VGND VPWR \$4438 \$4508 \$907 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$10990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$10992 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$10993 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$10994 VPWR \$4439 VPWR \$4671 VGND \$3993 \$2472 VGND sky130_fd_sc_hd__o21a_1
X$10995 VPWR \$4697 VGND VPWR \$4733 \$4726 \$1962 \$3833 VGND
+ sky130_fd_sc_hd__o22a_1
X$10996 VPWR VGND \$2336 VPWR \$3649 \$4697 VGND sky130_fd_sc_hd__nor2_2
X$10997 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$10998 VPWR \$4726 VGND \$3916 \$1998 VPWR VGND sky130_fd_sc_hd__or2_1
X$10999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11000 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11001 VPWR VPWR \$4733 VGND \$4726 \$4475 \$4445 VGND sky130_fd_sc_hd__o21ai_1
X$11002 VPWR VGND VPWR \$4652 \$4210 VGND sky130_fd_sc_hd__inv_2
X$11003 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11005 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11007 VPWR \$2741 VGND VPWR \$4210 \$4698 VGND sky130_fd_sc_hd__or2_4
X$11008 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11009 VPWR \$4139 VPWR VGND \$2742 \$4698 VGND sky130_fd_sc_hd__or2_2
X$11010 VPWR VGND VPWR \$4512 \$4698 VGND sky130_fd_sc_hd__inv_2
X$11011 VPWR \$4445 VPWR VGND \$4006 \$4698 VGND sky130_fd_sc_hd__or2_2
X$11012 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11013 VPWR VGND VPWR \$4412 \$3342 VGND sky130_fd_sc_hd__inv_2
X$11014 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11015 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11016 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11017 VGND \$4223 \$4757 \$4249 \$2700 \$4734 \$4604 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$11018 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11019 VPWR \$4712 VPWR VGND \$4578 \$4577 \$4252 VGND sky130_fd_sc_hd__or3_1
X$11020 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11021 VPWR \$4713 VGND \$4735 \$4712 VPWR VGND sky130_fd_sc_hd__or2_1
X$11022 VGND \$4674 \$4663 \$4664 \$4412 \$4713 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$11023 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11025 VPWR \$4672 VGND VPWR \$3342 \$4673 \$4673 \$1979 VGND
+ sky130_fd_sc_hd__o22a_1
X$11026 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11027 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11028 VPWR VGND \$4603 VPWR \$4736 \$4139 VGND sky130_fd_sc_hd__nor2_2
X$11029 VPWR VPWR \$4529 VGND \$4615 \$4664 \$4736 \$4699 VGND
+ sky130_fd_sc_hd__a211o_1
X$11030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11031 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11032 VPWR \$4672 VGND \$4688 VPWR \$4700 VGND sky130_fd_sc_hd__or2b_1
X$11033 VPWR \$4570 VGND \$1963 VPWR \$4623 VGND sky130_fd_sc_hd__nor2_1
X$11034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11036 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11037 VPWR \$4571 VGND \$4737 \$4738 VPWR VGND sky130_fd_sc_hd__or2_1
X$11038 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11039 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11040 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11041 VPWR \$4714 VGND \$4700 \$4699 VPWR VGND sky130_fd_sc_hd__or2_1
X$11042 VPWR \$4269 VPWR VGND \$4739 \$4676 \$4699 VGND sky130_fd_sc_hd__or3_1
X$11043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11044 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11045 VPWR \$4728 VPWR VGND \$4665 \$4727 \$4714 VGND sky130_fd_sc_hd__or3_1
X$11046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11048 VPWR \$4740 VGND VPWR \$4728 VGND sky130_fd_sc_hd__clkbuf_1
X$11049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11050 VGND \$3507 \$4741 \$4740 \$1724 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$11051 VPWR VPWR VGND \$3702 \$4715 VGND sky130_fd_sc_hd__clkbuf_2
X$11052 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11053 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11054 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11055 VPWR VGND \$4555 \$3732 \$4689 \$4716 \$4530 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11056 VGND \$2777 \$4689 \$4216 \$4716 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11057 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11058 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11060 VGND \$2777 \$4702 \$4216 \$4729 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11061 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11062 VPWR VGND \$4701 \$4023 \$4702 \$4729 \$4677 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11063 VPWR \$3883 \$4689 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11064 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11065 VPWR VGND VPWR \$2957 \$4702 VGND sky130_fd_sc_hd__inv_2
X$11066 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11067 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11069 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11070 VGND \$4353 \$4703 \$4406 \$4742 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11071 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11072 VPWR VPWR VGND \$4289 \$4717 VGND sky130_fd_sc_hd__clkbuf_2
X$11073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11074 VPWR VGND VPWR \$2597 \$4703 VGND sky130_fd_sc_hd__inv_2
X$11075 VGND \$4353 \$4704 \$4406 \$4743 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11076 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11077 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11079 VPWR VGND VPWR \$2539 \$4704 VGND sky130_fd_sc_hd__inv_2
X$11080 VGND \$4374 \$4406 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$11081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11082 VPWR VGND VPWR \$3017 \$4744 VGND sky130_fd_sc_hd__inv_2
X$11083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11085 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11086 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11087 VGND \$4353 \$4705 \$4406 \$4718 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11088 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11089 VPWR VGND \$4654 \$3711 \$4705 \$4718 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11090 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11091 VPWR VGND VPWR \$3265 \$4705 VGND sky130_fd_sc_hd__inv_2
X$11092 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11094 VGND \$4353 \$4690 \$4377 \$4719 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11095 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11096 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11097 VPWR VGND \$4654 \$1179 \$4690 \$4719 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11099 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11101 VPWR VGND VPWR \$2599 \$4690 VGND sky130_fd_sc_hd__inv_2
X$11102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11103 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11104 VPWR VGND \$4707 \$4023 \$4669 \$4668 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11105 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11106 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11107 VPWR \$2790 \$4745 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11108 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11109 VPWR \$4720 VGND \$2789 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$11110 VGND \$4353 \$4679 \$4377 \$4730 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11111 VPWR VGND \$4707 \$1594 \$4679 \$4730 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11112 VPWR VGND \$4706 VPWR \$4720 VGND sky130_fd_sc_hd__clkbuf_4
X$11113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11115 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11116 VGND \$4353 \$4680 \$4424 \$4691 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11118 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11119 VPWR VGND \$4681 \$1594 \$4683 \$4721 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11120 VGND \$4353 \$4683 \$4424 \$4721 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11121 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11123 VGND \$4353 \$4684 \$4424 \$4722 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11124 VPWR VGND \$4681 \$1179 \$4684 \$4722 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11125 VPWR VGND \$4682 VPWR \$4692 VGND sky130_fd_sc_hd__clkbuf_4
X$11126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11128 VPWR \$3715 \$4746 VPWR \$4670 VGND \$1125 \$3869 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$11129 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11132 VPWR VGND \$4707 \$184 \$4747 \$4748 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11134 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11137 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11140 VPWR \$4693 VGND \$2667 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$11141 VPWR VGND VPWR \$3927 \$4747 VGND sky130_fd_sc_hd__inv_2
X$11142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11143 VPWR \$4694 VGND VPWR \$3927 \$2789 \$4628 \$2447 VGND
+ sky130_fd_sc_hd__o22a_1
X$11144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11146 VGND \$4280 \$4694 \$3480 \$2751 \$2918 \$4030 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11148 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11150 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11151 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11152 VPWR \$3168 \$4756 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11153 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11154 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11156 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11157 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11158 VPWR VGND VPWR \$4146 \$4708 VGND sky130_fd_sc_hd__inv_2
X$11159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11162 VPWR VGND \$4709 \$184 \$4708 \$4723 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11163 VGND \$2989 \$4708 \$4427 \$4723 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11166 VPWR VGND \$4709 \$1179 \$4649 \$4685 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11167 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11169 VPWR VGND \$4709 \$354 \$4613 \$4658 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11172 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11174 VPWR \$1588 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11176 VPWR \$4749 VGND \$2117 \$2474 VPWR VGND sky130_fd_sc_hd__or2_1
X$11177 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11178 VPWR \$1588 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11179 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11180 VGND \$4724 \$345 \$4695 \$4239 \$2474 VPWR VPWR VGND
+ sky130_fd_sc_hd__a211o_4
X$11181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11183 VGND \$4695 \$3611 \$3924 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$11184 VPWR \$2869 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11185 VGND \$4731 \$2869 \$4751 \$4750 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$11186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11187 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11188 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11190 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11191 VGND \$4731 \$2863 mgmt_gpio_out[13] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$11192 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11195 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11199 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11201 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11202 VPWR VGND wb_dat_o[5] VPWR \$4175 VGND sky130_fd_sc_hd__buf_2
X$11203 VGND \$4175 \$3277 \$4192 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$11204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11206 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11207 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11209 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11210 VGND \$4194 \$4210 \$4211 \$4149 \$3916 \$1963 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$11211 VPWR \$4149 VGND \$3057 \$2996 VPWR VGND sky130_fd_sc_hd__or2_1
X$11212 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11213 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11214 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11215 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11216 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11217 VPWR \$4177 VGND \$4212 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$11218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11220 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11221 VGND \$4213 \$4249 \$4061 \$2815 \$4210 \$4212 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$11222 VPWR \$4214 VGND \$4213 \$3502 VPWR \$3995 VGND sky130_fd_sc_hd__o21ai_2
X$11223 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11225 VPWR \$4062 VGND \$4214 \$4249 VPWR VGND sky130_fd_sc_hd__or2_1
X$11226 VPWR \$4077 VGND \$4214 \$4250 VPWR VGND sky130_fd_sc_hd__or2_1
X$11227 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11228 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11231 VPWR \$4251 VGND \$4078 \$4250 VPWR VGND sky130_fd_sc_hd__or2_1
X$11232 VPWR \$4178 VGND \$4195 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$11233 VPWR \$4215 VGND \$2700 \$4251 VPWR VGND sky130_fd_sc_hd__or2_1
X$11234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11235 VPWR \$4179 VGND \$2741 \$4251 VPWR VGND sky130_fd_sc_hd__or2_1
X$11236 VPWR VPWR \$3709 VGND \$4195 \$4252 \$3454 VGND sky130_fd_sc_hd__o21ai_1
X$11237 VPWR \$4180 VGND \$4151 \$4215 VPWR VGND sky130_fd_sc_hd__or2_1
X$11238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11239 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11240 VPWR \$5004 VGND \$4196 \$4152 VPWR VGND sky130_fd_sc_hd__or2_1
X$11241 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11242 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11243 VPWR VPWR \$4179 VGND \$4151 \$4140 \$4180 VGND sky130_fd_sc_hd__o21ai_1
X$11244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11246 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11249 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11251 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11252 VGND \$2777 \$4254 \$4216 \$4233 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11254 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11255 VGND \$2777 \$4198 \$4216 \$4217 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11256 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11257 VPWR VGND \$4234 \$3694 \$4198 \$4217 \$4224 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11260 VPWR \$4199 VGND \$3703 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$11261 VPWR VPWR VGND \$4199 \$4224 VGND sky130_fd_sc_hd__clkbuf_2
X$11262 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11263 VPWR \$4255 VGND \$3562 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$11264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11266 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11268 VPWR VGND \$4183 \$3732 \$4171 \$4182 \$4185 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11269 VGND \$2777 \$4184 \$3921 \$4200 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11271 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11272 VPWR VPWR VGND \$4201 \$4185 VGND sky130_fd_sc_hd__clkbuf_2
X$11273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11275 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11276 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11280 VGND \$2777 \$4202 \$3921 \$4225 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11281 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11282 VPWR \$4225 VGND VPWR \$4218 VGND sky130_fd_sc_hd__clkbuf_1
X$11283 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11284 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11285 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11287 VPWR \$1333 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11288 VGND \$1341 \$1333 \$4226 \$4202 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$11289 VPWR \$4186 VPWR VGND \$1571 \$1425 \$345 VGND sky130_fd_sc_hd__or3_1
X$11290 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11291 VPWR VGND VPWR \$4235 \$4202 VGND sky130_fd_sc_hd__inv_2
X$11292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11293 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11294 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11295 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11296 VPWR \$4256 VGND VPWR \$2783 \$3556 \$2840 \$3271 VGND
+ sky130_fd_sc_hd__o22a_1
X$11297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11299 VPWR \$4228 VGND VPWR \$4117 \$2229 \$3395 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$11300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11301 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11302 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11303 VGND \$4227 \$1571 \$1425 \$4235 \$2474 \$4236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$11304 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11305 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11306 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11307 VGND \$4229 \$4227 \$4237 \$2614 \$3042 \$3551 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11308 VPWR VGND VPWR \$3577 \$4219 \$4313 \$4203 \$3764 VGND
+ sky130_fd_sc_hd__and4_1
X$11309 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11310 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11311 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11312 VPWR VGND VPWR \$4219 \$4220 \$4204 \$3205 \$4229 VGND
+ sky130_fd_sc_hd__and4_1
X$11313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11314 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11315 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11317 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11318 VPWR \$4238 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11319 VGND \$4220 \$4238 \$4230 \$4239 \$2918 \$4119 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11322 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11323 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11324 VGND \$4221 \$4240 \$4134 \$2525 \$2458 \$4241 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11325 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11328 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11329 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11330 VGND \$4231 \$4242 \$4028 \$1065 \$880 \$4107 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11333 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11335 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11336 VGND \$4222 \$4228 \$3447 \$2330 \$2219 \$3673 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11337 VPWR VGND VPWR \$4206 \$4205 \$4222 \$4231 \$3238 VGND
+ sky130_fd_sc_hd__and4_1
X$11338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11341 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11344 VPWR \$4259 VGND VPWR \$4258 \$2456 \$4243 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$11345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11347 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11348 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11350 VPWR \$4207 VGND VPWR \$1077 \$2135 \$3254 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$11351 VPWR \$4208 VGND VPWR \$1812 \$2456 \$4146 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$11352 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11354 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11355 VPWR \$4260 VGND VPWR \$2629 \$2456 \$4244 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$11356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11358 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11363 VPWR VGND VPWR \$4031 \$4245 VGND sky130_fd_sc_hd__inv_2
X$11364 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11366 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11367 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11369 VPWR VGND VPWR \$3209 \$3609 VGND sky130_fd_sc_hd__inv_4
X$11370 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11372 VPWR \$4261 VPWR VGND \$3209 \$464 VGND sky130_fd_sc_hd__or2_2
X$11373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11375 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11380 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11381 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11382 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11383 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11384 VPWR \$3748 \$4246 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11389 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11390 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11391 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11392 VPWR \$3929 \$4247 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11394 VGND \$2989 \$4247 \$4165 \$4262 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11395 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11400 VPWR VGND \$4248 \$2897 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$11401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11404 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11405 VGND \$1830 \$1860 \$1376 \$1827 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$11406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11407 VPWR \$1875 \$1885 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11408 VPWR \$1885 VGND VPWR sram_ro_data[22] VGND sky130_fd_sc_hd__clkbuf_1
X$11409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11410 VPWR VGND \$1514 \$1806 \$1860 \$1827 \$1473 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11412 VPWR \$1830 VGND VPWR \$1828 VGND sky130_fd_sc_hd__clkbuf_1
X$11413 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11414 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11418 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11419 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11420 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11421 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11426 VPWR \$1900 VGND \$1886 \$1898 VPWR VGND sky130_fd_sc_hd__or2_1
X$11427 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11428 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11429 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11431 VPWR \$1901 VGND \$1887 \$1900 VPWR VGND sky130_fd_sc_hd__or2_1
X$11432 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11433 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11436 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11438 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11439 VPWR VGND \$1725 \$1550 \$1850 \$1832 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11440 VPWR VGND \$1725 \$1488 \$1888 \$1849 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11444 VPWR VPWR VGND \$1902 \$381 VGND sky130_fd_sc_hd__clkbuf_2
X$11445 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11447 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11449 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11451 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11453 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11454 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11458 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11459 VPWR VGND \$1752 \$281 \$1905 \$1904 \$1774 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11462 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11463 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11464 VPWR VGND VPWR \$1851 \$1773 VGND sky130_fd_sc_hd__inv_2
X$11465 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11466 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11467 VPWR \$1862 VGND VPWR \$1852 \$1729 \$1851 \$1713 VGND
+ sky130_fd_sc_hd__o22a_1
X$11468 VGND \$1876 \$1862 \$709 \$927 \$1297 \$1805 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11469 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11470 VGND \$856 \$1835 \$1861 \$1834 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11471 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11472 VPWR \$1906 VGND \$1444 \$1571 VPWR VGND sky130_fd_sc_hd__or2_1
X$11473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11476 VPWR VGND \$1567 \$183 \$1889 \$1877 \$1568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11477 VGND \$856 \$1889 \$1863 \$1877 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11478 VPWR VGND VPWR \$1907 \$1835 VGND sky130_fd_sc_hd__inv_2
X$11479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11480 VPWR VGND VPWR \$1853 \$1889 VGND sky130_fd_sc_hd__inv_2
X$11481 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11483 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11484 VPWR \$1342 VGND VPWR \$1810 \$1059 VGND sky130_fd_sc_hd__or2_4
X$11485 VPWR \$1908 VGND VPWR \$1611 \$1776 \$1076 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$11486 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11487 VPWR \$1864 VGND VPWR \$1807 \$1776 \$1004 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$11488 VGND \$1908 \$1569 \$1715 \$1754 \$1259 \$1878 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$11489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11492 VGND \$1866 \$1789 \$1853 \$1715 \$1754 \$1236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11493 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11495 VPWR \$1865 VGND VPWR \$726 \$1060 \$1853 \$1613 VGND
+ sky130_fd_sc_hd__o22a_1
X$11496 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11497 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11498 VPWR \$1490 VGND VPWR \$1890 \$1356 VGND sky130_fd_sc_hd__or2_4
X$11499 VPWR \$1490 VGND VPWR \$1867 \$1283 VGND sky130_fd_sc_hd__or2_4
X$11500 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11502 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11503 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11504 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11505 VGND \$1844 \$1402 \$1875 \$1554 \$1879 \$1880 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11507 VPWR \$1598 VGND VPWR \$1845 \$1283 VGND sky130_fd_sc_hd__or2_4
X$11508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11509 VPWR \$1490 VGND VPWR \$1879 \$1329 VGND sky130_fd_sc_hd__or2_4
X$11510 VPWR \$1490 VGND VPWR \$1839 \$1258 VGND sky130_fd_sc_hd__or2_4
X$11511 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11513 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11516 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11517 VGND \$1777 \$1891 \$1892 \$1645 \$1643 \$1807 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11518 VGND \$1868 \$1840 \$1854 \$1841 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$11519 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11520 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11521 VPWR \$1909 VGND VPWR \$1807 \$1793 \$1869 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$11522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11524 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11526 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11528 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11529 VPWR VGND \$1572 \$200 \$1910 \$1926 \$1592 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11530 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11532 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11533 VPWR VPWR VGND \$1911 \$1592 VGND sky130_fd_sc_hd__clkbuf_2
X$11534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11535 VGND \$358 \$1627 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$11536 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11537 VPWR VGND VPWR \$1869 \$1796 VGND sky130_fd_sc_hd__inv_2
X$11538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11539 VGND \$1854 \$1846 \$335 \$456 \$1819 \$1855 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11540 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11541 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11542 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11544 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11545 VPWR \$1881 VGND VPWR \$977 \$1114 \$1802 \$2180 VGND
+ sky130_fd_sc_hd__o22a_1
X$11546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11547 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11548 VGND \$1912 \$1881 \$871 \$848 \$1676 \$1893 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11549 VGND \$1870 \$1822 \$1606 \$520 \$1839 \$1856 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11552 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11553 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11554 VPWR \$1871 VGND \$1779 \$1766 VPWR VGND sky130_fd_sc_hd__or2_1
X$11555 VGND \$1871 \$1954 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$11556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11558 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11559 VPWR \$1913 VPWR VGND \$1128 \$1882 \$1705 VGND sky130_fd_sc_hd__or3_1
X$11560 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11561 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11563 VPWR \$1825 VPWR VGND \$1798 \$1746 \$1766 VGND sky130_fd_sc_hd__or3_1
X$11564 VGND \$1799 \$1955 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$11565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11566 VGND \$1894 \$1914 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$11567 VPWR \$1894 VGND \$1779 \$1782 VPWR VGND sky130_fd_sc_hd__or2_1
X$11568 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11569 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11572 VGND \$1152 \$1662 \$541 \$1800 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_2
X$11573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11577 VGND \$516 \$1857 \$1273 \$1872 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11578 VPWR VGND \$1680 \$386 \$1857 \$1872 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11580 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11581 VPWR VGND \$1680 \$1594 \$1858 \$1873 \$1681 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11582 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11583 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11584 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11585 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11586 VGND \$516 \$1858 \$1273 \$1873 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11588 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11590 VPWR VGND \$1311 \$354 \$1848 \$1826 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11591 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11592 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11594 VGND \$1884 \$354 \$1848 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$11595 VGND \$358 \$1874 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$11596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11597 VPWR \$1916 VGND VPWR \$1884 \$1363 \$1895 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$11598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11599 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11600 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11606 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11607 VPWR \$1564 VGND VPWR sram_ro_data[18] VGND sky130_fd_sc_hd__clkbuf_1
X$11608 VPWR \$1577 VGND VPWR sram_ro_data[17] VGND sky130_fd_sc_hd__clkbuf_1
X$11609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11611 VPWR \$1632 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$11612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11613 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11615 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11616 VGND \$1596 \$1633 \$381 \$1618 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$11617 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11619 VPWR \$1578 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$11620 VPWR \$1596 VGND VPWR \$1578 VGND sky130_fd_sc_hd__clkbuf_1
X$11621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11622 VGND \$1524 \$1619 \$1633 \$1186 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$11623 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11624 VGND \$1579 \$1580 \$1376 \$1597 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$11625 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11628 VPWR VGND \$1053 \$1581 \$1580 \$1597 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11629 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11630 VGND \$1634 \$1583 \$1580 \$1620 \$1609 \$1610 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$11631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11633 VPWR \$1583 VPWR \$1582 VGND \$1610 \$1580 VGND sky130_fd_sc_hd__o21a_1
X$11634 VPWR \$1610 VPWR VGND \$1580 \$1583 VGND sky130_fd_sc_hd__nand2_1
X$11635 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11636 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11639 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11640 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11642 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11646 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11647 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11648 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11649 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11650 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11651 VPWR VGND \$1399 \$281 \$1540 \$1539 \$1417 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11652 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11653 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11654 VGND \$856 \$1566 \$1370 \$1552 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11655 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11656 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11657 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11658 VPWR \$1611 \$1527 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11659 VPWR VPWR VGND \$1621 \$1417 VGND sky130_fd_sc_hd__clkbuf_2
X$11660 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11661 VPWR \$1637 \$1566 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11665 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11668 VGND \$1506 \$1598 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$11669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11671 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11672 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11673 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11674 VPWR VGND VPWR \$1567 \$1568 VGND sky130_fd_sc_hd__inv_2
X$11675 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11677 VPWR VGND \$1567 \$293 \$1622 \$1638 \$1568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11678 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11679 VPWR \$1623 VGND \$1613 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$11680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11681 VPWR VPWR VGND \$1623 \$1568 VGND sky130_fd_sc_hd__clkbuf_2
X$11682 VPWR \$1613 VPWR VGND \$1401 \$1571 VGND sky130_fd_sc_hd__or2_2
X$11683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11684 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11685 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11686 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11687 VPWR \$1059 VGND VPWR \$1588 \$1248 VGND sky130_fd_sc_hd__or2_4
X$11688 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11689 VPWR \$1598 VGND VPWR \$1116 \$1434 VGND sky130_fd_sc_hd__or2_4
X$11690 VGND \$517 \$1569 \$1613 \$1116 \$1259 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$11691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11692 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11693 VPWR \$1599 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11694 VPWR \$1589 VGND VPWR \$1496 \$1297 \$1599 \$1588 VGND
+ sky130_fd_sc_hd__o22a_1
X$11695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11696 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11697 VGND \$1669 \$1589 \$1548 \$1554 \$744 \$770 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11699 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11700 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11701 VPWR \$1612 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11702 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11703 VPWR \$1600 VGND VPWR \$678 \$1114 \$1612 \$1125 VGND
+ sky130_fd_sc_hd__o22a_1
X$11704 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11705 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11706 VPWR \$1612 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11707 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11708 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11709 VPWR \$1624 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11710 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11711 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11712 VGND \$1640 \$1381 \$899 \$1238 \$1624 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$11713 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11714 VPWR \$1598 VGND VPWR \$1625 \$1445 VGND sky130_fd_sc_hd__or2_4
X$11715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11718 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11722 VGND \$1585 \$1601 \$1625 \$286 \$420 \$1590 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_4
X$11723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11726 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11729 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11730 VPWR VGND \$1572 \$1179 \$1591 \$1573 \$1592 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11731 VPWR \$1602 \$1591 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11732 VPWR VGND \$1572 \$294 \$1626 \$1614 \$1592 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11733 VPWR VGND VPWR \$1572 \$1592 VGND sky130_fd_sc_hd__inv_2
X$11734 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11736 VGND \$1152 \$1626 \$1627 \$1614 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11740 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11741 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11744 VPWR VGND VPWR \$1603 \$1530 VGND sky130_fd_sc_hd__inv_2
X$11745 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11746 VGND \$1152 \$1604 \$1203 \$1586 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11748 VPWR VGND VPWR \$1628 \$1604 VGND sky130_fd_sc_hd__inv_2
X$11749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11750 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11751 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11752 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11753 VGND \$1152 \$1593 \$1203 \$1605 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11754 VPWR VGND \$1170 \$411 \$1593 \$1605 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11755 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11757 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11758 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11759 VPWR VGND VPWR \$2630 \$1519 VGND sky130_fd_sc_hd__inv_2
X$11760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11762 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11763 VGND \$1629 \$1011 \$1798 \$1673 \$1205 \$1630 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$11764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11767 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11770 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11771 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11772 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11773 VPWR \$1631 VGND \$1575 \$1576 VPWR VGND sky130_fd_sc_hd__or2_1
X$11774 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11775 VPWR \$1546 VGND VPWR \$1780 \$1534 VGND sky130_fd_sc_hd__or2_4
X$11776 VPWR \$1784 VGND \$1546 \$1576 VPWR VGND sky130_fd_sc_hd__or2_1
X$11777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11778 VPWR VGND VPWR \$1575 \$1546 VGND sky130_fd_sc_hd__inv_2
X$11779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11781 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11782 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11783 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11784 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11785 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11786 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11788 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11789 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11791 VPWR VGND \$1311 \$1594 \$1595 \$1607 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11792 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11793 VGND \$516 \$1595 \$1273 \$1607 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11794 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11795 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11796 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11797 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11799 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11800 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11801 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11803 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11804 VGND \$4264 \$3277 \$4324 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$11805 VPWR VGND wb_dat_o[7] VPWR \$4349 VGND sky130_fd_sc_hd__buf_2
X$11806 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11807 VGND \$4349 \$3277 \$4366 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$11808 VPWR \$4366 VGND VPWR \$4349 \$3531 \$1619 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$11809 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11810 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11811 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11812 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11813 VGND \$4367 \$3742 \$3332 \$3805 \$4350 \$2552 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_4
X$11814 VPWR VGND \$4351 \$4359 \$4325 VPWR \$4034 \$4350 VGND
+ sky130_fd_sc_hd__or4b_2
X$11815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11817 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11818 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11819 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11820 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11821 VPWR \$3484 \$4396 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11824 VPWR \$4337 VGND \$4151 VPWR \$4210 VGND sky130_fd_sc_hd__nor2_1
X$11825 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11826 VPWR \$3249 VGND \$4050 \$4368 VPWR VGND sky130_fd_sc_hd__or2_1
X$11827 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11828 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11829 VPWR \$4352 VGND \$4368 \$4078 VPWR VGND sky130_fd_sc_hd__or2_1
X$11830 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11831 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11833 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11834 VPWR VPWR VGND \$3702 \$4266 VGND sky130_fd_sc_hd__clkbuf_2
X$11835 VPWR VGND \$3710 VPWR \$4352 VGND sky130_fd_sc_hd__buf_2
X$11836 VGND \$4369 \$4397 \$3484 \$3858 \$3860 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$11837 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11839 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11840 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11842 VPWR \$4371 VGND \$3710 \$2700 VPWR VGND sky130_fd_sc_hd__or2_1
X$11843 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11844 VPWR \$4372 VGND \$4370 \$4197 VPWR VGND sky130_fd_sc_hd__or2_1
X$11845 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11846 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11847 VPWR \$4373 VGND \$4372 \$4286 VPWR VGND sky130_fd_sc_hd__or2_1
X$11848 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11849 VPWR \$4286 VGND \$4310 VPWR \$2700 VGND sky130_fd_sc_hd__nor2_1
X$11850 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11852 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11853 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11855 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11857 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11858 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11859 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11860 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11862 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11863 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11864 VPWR VGND VPWR \$4234 \$4224 VGND sky130_fd_sc_hd__inv_2
X$11865 VGND \$2777 \$4327 \$3921 \$4328 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11866 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11867 VPWR \$3840 \$4382 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$11868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11870 VGND \$4353 \$4354 \$3921 \$4360 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11871 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11872 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11873 VGND \$2777 \$4353 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$11874 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11875 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11876 VPWR VGND VPWR \$2971 \$4354 VGND sky130_fd_sc_hd__inv_2
X$11877 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11879 VGND \$4374 \$3921 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$11880 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11884 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11887 VPWR \$4375 VGND \$1810 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$11888 VPWR VPWR VGND \$4375 \$4376 VGND sky130_fd_sc_hd__clkbuf_2
X$11889 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11890 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11891 VPWR VGND \$4405 \$4023 \$4361 \$4355 \$4376 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11892 VGND \$4353 \$4361 \$3921 \$4355 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11893 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11894 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11895 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11896 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11897 VPWR VGND VPWR \$1837 \$4361 VGND sky130_fd_sc_hd__inv_2
X$11898 VPWR VGND VPWR \$3935 \$4384 VGND sky130_fd_sc_hd__inv_2
X$11899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11900 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11901 VPWR \$4338 VGND \$1819 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$11902 VGND \$4353 \$4386 \$4377 \$4362 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11903 VPWR VGND \$4363 VPWR \$4338 VGND sky130_fd_sc_hd__clkbuf_4
X$11904 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11905 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11908 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11909 VPWR \$4339 VGND VPWR \$4275 \$2135 \$2804 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$11910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11911 VGND \$4340 \$4339 \$4119 \$1065 \$880 \$3161 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11912 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11913 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11915 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11916 VPWR VGND VPWR \$4276 \$4330 \$4341 \$4340 \$3671 VGND
+ sky130_fd_sc_hd__and4_1
X$11917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11921 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11922 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11927 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11928 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11929 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11930 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11932 VGND \$4353 \$4389 \$4424 \$4378 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11933 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11934 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11935 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11937 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11938 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11939 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11940 VPWR VGND VPWR \$4343 \$4333 \$4342 \$4332 \$3109 VGND
+ sky130_fd_sc_hd__and4_1
X$11941 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11942 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$11943 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11944 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11945 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11946 VPWR \$4344 VGND VPWR \$4294 \$2135 \$3404 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$11947 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11949 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11950 VGND \$4345 \$4344 \$3629 \$1065 \$880 \$3587 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$11951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11952 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11953 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11954 VPWR VGND VPWR \$4364 \$4334 \$4356 \$4345 \$3646 VGND
+ sky130_fd_sc_hd__and4_1
X$11955 VPWR \$691 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$11956 VGND \$3736 \$4364 \$4454 VPWR \$691 VPWR VGND sky130_fd_sc_hd__nand3_4
X$11957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11959 VPWR VGND \$4358 VPWR \$4335 VGND sky130_fd_sc_hd__buf_2
X$11960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11961 VPWR VGND \$4357 \$184 \$4245 \$4297 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11963 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11964 VPWR VGND \$4357 \$1594 \$4189 \$4346 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11965 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11966 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$11969 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11971 VGND \$2989 \$4282 \$4427 \$4336 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$11972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11975 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11976 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11977 VPWR VGND \$4303 \$1179 \$4246 \$4322 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11978 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11980 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11982 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$11983 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11984 VGND \$2989 \$4347 \$4165 \$4365 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$11985 VPWR VGND VPWR \$3581 \$4347 VGND sky130_fd_sc_hd__inv_2
X$11986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11987 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11988 VPWR VGND \$3872 \$1171 \$4347 \$4365 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$11989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$11990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$11991 VGND \$2989 \$4285 \$4165 \$4348 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$11992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11993 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$11994 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11995 VPWR \$4379 VGND VPWR \$4380 VGND sky130_fd_sc_hd__clkbuf_1
X$11996 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$11997 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11998 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$11999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12001 VGND \$4538 \$4651 \$4643 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$12002 VPWR VGND wb_dat_o[14] VPWR \$4950 VGND sky130_fd_sc_hd__buf_2
X$12003 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12004 VPWR \$4643 VGND VPWR \$4538 \$4508 \$2057 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$12005 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12006 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12007 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12008 VPWR \$3854 VPWR VGND \$4671 \$4474 VGND sky130_fd_sc_hd__or2_2
X$12009 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12011 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12012 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12013 VPWR \$4474 VGND \$4644 \$4359 VPWR \$4632 VGND sky130_fd_sc_hd__o21ai_2
X$12014 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12015 VPWR \$4644 VGND \$4615 VPWR \$4645 VGND sky130_fd_sc_hd__nor2_1
X$12016 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12018 VGND \$4549 \$4511 \$4726 \$4645 VPWR VPWR \$4652 VGND
+ sky130_fd_sc_hd__or4bb_1
X$12019 VPWR \$4652 VGND \$4633 \$4350 VPWR \$4646 VGND sky130_fd_sc_hd__o21ai_2
X$12020 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12021 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12023 VGND \$4687 \$4652 \$4645 \$4662 \$4308 VPWR VPWR VGND
+ sky130_fd_sc_hd__o31a_1
X$12024 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12025 VPWR VGND VPWR \$4645 \$4445 VGND sky130_fd_sc_hd__inv_2
X$12026 VPWR \$4306 VGND \$4615 VPWR \$4662 VGND sky130_fd_sc_hd__nor2_1
X$12027 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12028 VPWR VGND VPWR \$4662 \$4139 VGND sky130_fd_sc_hd__inv_2
X$12029 VPWR VPWR \$4210 VGND \$4151 \$4308 \$4214 VGND sky130_fd_sc_hd__o21ai_1
X$12030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12031 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12032 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12033 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12034 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12036 VPWR \$3857 \$4663 \$4646 VGND VPWR \$3343 VGND sky130_fd_sc_hd__and3_2
X$12037 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12038 VPWR VGND VPWR \$4604 \$4370 VGND sky130_fd_sc_hd__inv_2
X$12039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12040 VPWR \$4412 \$4664 \$4512 VGND VPWR \$4665 VGND sky130_fd_sc_hd__and3_2
X$12041 VPWR \$4550 \$4672 VPWR \$4603 \$4445 \$1962 VGND \$4673 VGND
+ sky130_fd_sc_hd__o221ai_1
X$12042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12043 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12044 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12046 VPWR \$4688 VPWR VGND \$4267 \$4153 \$4674 VGND sky130_fd_sc_hd__or3_1
X$12047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12048 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12049 VPWR \$4552 VGND \$1998 VPWR \$4623 VGND sky130_fd_sc_hd__nor2_1
X$12050 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12051 VPWR \$4520 \$4589 \$4571 VPWR VGND \$4675 \$4503 VGND
+ sky130_fd_sc_hd__or4_1
X$12052 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12054 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12055 VPWR \$4666 \$4553 VGND \$4699 VPWR \$4312 \$4519 VGND
+ sky130_fd_sc_hd__or4_2
X$12056 VPWR \$4666 VPWR VGND \$4552 \$4738 \$4676 VGND sky130_fd_sc_hd__or3_1
X$12057 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12058 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12059 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12060 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12061 VGND \$2777 \$4634 \$4216 \$4647 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12062 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12063 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12065 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12066 VPWR VGND VPWR \$3910 \$4634 VGND sky130_fd_sc_hd__inv_2
X$12067 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12069 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12071 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12072 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12073 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12074 VPWR VPWR VGND \$4635 \$4677 VGND sky130_fd_sc_hd__clkbuf_2
X$12075 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12076 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12077 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12078 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12079 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12084 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12085 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12087 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12088 VPWR \$4678 VPWR VGND \$3553 \$345 VGND sky130_fd_sc_hd__or2_2
X$12089 VPWR VPWR VGND \$4637 \$4782 VGND sky130_fd_sc_hd__clkbuf_2
X$12090 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12092 VGND \$4353 \$4624 \$4406 \$4653 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12093 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12095 VPWR VGND \$4654 \$3732 \$4624 \$4653 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12096 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12097 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12098 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12099 VPWR VGND \$4667 VPWR \$4638 VGND sky130_fd_sc_hd__buf_2
X$12100 VPWR VGND \$4654 \$411 \$4648 \$4655 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12102 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12103 VGND \$4353 \$4648 \$4377 \$4655 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12105 VGND \$4353 \$4669 \$4377 \$4668 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12106 VGND \$4374 \$4377 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12107 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12108 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12111 VPWR \$2752 \$4679 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12112 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12114 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12115 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12116 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12117 VPWR VGND \$4680 \$1730 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$12118 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12119 VPWR VGND \$4681 \$4023 \$4680 \$4691 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12120 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12122 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12123 VPWR VGND VPWR \$2561 \$4683 VGND sky130_fd_sc_hd__inv_2
X$12124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12125 VPWR \$3540 \$4684 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12126 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12127 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12128 VPWR \$4692 VGND \$1676 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$12129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12131 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12132 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12134 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12135 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12136 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12137 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12138 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12139 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12142 VPWR \$4525 VGND VPWR \$3544 \$1561 \$4627 \$2667 VGND
+ sky130_fd_sc_hd__o22a_1
X$12143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12146 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12147 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12150 VGND \$4353 \$4610 \$4427 \$4656 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12151 VPWR VGND \$4357 \$1179 \$4610 \$4656 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12153 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12154 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12156 VPWR \$4657 VGND \$2986 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$12157 VPWR VGND \$4710 VPWR \$4657 VGND sky130_fd_sc_hd__clkbuf_4
X$12158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12159 VGND \$3952 \$4427 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12160 VGND \$1406 \$345 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$12161 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12162 VGND \$2989 \$4649 \$4165 \$4685 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12163 VPWR VGND VPWR \$4145 \$4649 VGND sky130_fd_sc_hd__inv_2
X$12164 VGND \$2989 \$4613 \$4165 \$4658 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12165 VPWR \$4686 VPWR VGND \$1588 \$345 VGND sky130_fd_sc_hd__or2_2
X$12166 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12167 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12168 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12169 VGND \$3924 \$2474 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$12170 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12171 VGND \$4629 \$3611 \$3869 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$12172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12173 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12174 VPWR VGND \$4659 VPWR \$4588 VGND sky130_fd_sc_hd__clkbuf_4
X$12175 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12176 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12177 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12178 VPWR VGND \$4650 \$1171 \$4564 \$4640 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12180 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12181 VPWR VGND \$4650 \$542 \$4641 \$4660 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12182 VGND \$2989 \$4641 \$4165 \$4660 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12184 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12185 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12187 VPWR \$4631 VGND VPWR \$2863 VGND sky130_fd_sc_hd__clkbuf_1
X$12188 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12192 VPWR \$2291 VGND VPWR sram_ro_data[28] VGND sky130_fd_sc_hd__clkbuf_1
X$12193 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12194 VPWR VGND VPWR \$1559 \$2319 VGND sky130_fd_sc_hd__inv_2
X$12195 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12196 VPWR VGND VPWR \$2310 \$2291 VGND sky130_fd_sc_hd__inv_2
X$12197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12200 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12201 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12206 VPWR \$2311 VGND \$2320 VPWR \$1999 VGND sky130_fd_sc_hd__nor2_1
X$12207 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12208 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12209 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12212 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12213 VPWR \$1887 VGND \$2320 VPWR \$2002 VGND sky130_fd_sc_hd__nor2_1
X$12214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12216 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12217 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12219 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12220 VPWR \$2312 VGND \$2337 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$12221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12222 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12223 VGND \$2026 \$2312 VPWR VPWR VGND sky130_fd_sc_hd__dlymetal6s2s_1
X$12224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12227 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12228 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12231 VGND \$856 \$2338 \$1750 \$2313 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12232 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12233 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12234 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12235 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12236 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12237 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12238 VPWR \$2292 \$2199 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12240 VGND \$856 \$2294 \$1370 \$2293 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12241 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12242 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12243 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12244 VPWR VGND \$2321 \$200 \$2294 \$2293 \$2322 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12246 VPWR VGND \$2321 \$293 \$2339 \$2340 \$2322 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12248 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12249 VPWR VGND VPWR \$2060 \$2294 VGND sky130_fd_sc_hd__inv_2
X$12250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12251 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12252 VGND \$463 \$1861 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12253 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12254 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12255 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12256 VGND \$856 \$2263 \$1861 \$2262 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12257 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12258 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12259 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12260 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12261 VPWR \$1435 VGND VPWR \$2314 \$1598 VGND sky130_fd_sc_hd__or2_4
X$12262 VPWR \$2247 \$2263 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12263 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12264 VGND \$2265 \$2279 \$988 \$2330 \$2219 \$2341 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12265 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12266 VGND \$2266 \$2264 \$2296 \$1065 \$880 \$2297 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12268 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12269 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12270 VGND \$2269 \$2280 \$725 \$785 \$2220 \$1950 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12272 VGND \$2267 \$2299 \$1081 \$2073 \$2096 \$2281 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12273 VPWR \$2315 VGND VPWR \$2225 \$1713 \$2342 \$2314 VGND
+ sky130_fd_sc_hd__o22a_1
X$12274 VPWR \$2343 VGND VPWR \$924 \$2724 \$2323 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$12275 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12276 VPWR \$2295 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12277 VPWR VGND VPWR \$2248 \$1716 \$2283 \$2282 \$2295 VGND
+ sky130_fd_sc_hd__and4_1
X$12278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12279 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12280 VPWR \$2344 VGND VPWR \$1236 \$2724 \$2383 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$12281 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12282 VGND \$2282 \$2284 \$2298 \$2043 \$1914 \$1019 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12283 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12284 VPWR \$2284 VGND VPWR \$2247 \$1966 \$2225 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$12285 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12286 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12287 VGND \$2317 \$2315 \$924 \$1116 \$859 \$1030 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12288 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12289 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12290 VGND \$2300 \$2239 \$770 \$1953 \$1987 \$1284 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12291 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12292 VPWR \$2345 VGND VPWR \$2324 \$2325 \$1349 \$1297 VGND
+ sky130_fd_sc_hd__o22a_1
X$12293 VPWR \$2299 VGND VPWR \$770 \$2045 \$1239 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$12294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12295 VPWR \$1598 VGND VPWR \$2162 \$1258 VGND sky130_fd_sc_hd__or2_4
X$12296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12297 VGND \$2301 \$2270 \$687 \$1953 \$1987 \$920 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12299 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12300 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12301 VPWR VPWR VGND \$2346 \$1446 VGND sky130_fd_sc_hd__clkbuf_2
X$12302 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12304 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12305 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12306 VGND \$2318 \$2326 \$2285 \$2065 \$2046 \$1239 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12307 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12308 VPWR \$2302 VGND VPWR \$1284 \$1956 \$1602 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$12309 VPWR \$2326 VGND VPWR \$1419 \$1793 \$1602 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$12310 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12311 VGND \$2228 \$2302 \$2285 \$2047 \$2048 \$756 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12312 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12313 VGND \$2328 \$2250 \$2327 \$2047 \$2048 \$796 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12316 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12317 VPWR \$2303 VGND VPWR \$1778 \$1890 \$1943 \$2180 VGND
+ sky130_fd_sc_hd__o22a_1
X$12318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12319 VPWR VGND VPWR \$2327 \$2329 VGND sky130_fd_sc_hd__inv_2
X$12320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12321 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12322 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12323 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12324 VPWR \$2304 VGND VPWR \$2286 \$1561 \$1701 \$848 VGND
+ sky130_fd_sc_hd__o22a_1
X$12325 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12326 VPWR VGND VPWR \$2285 \$2305 VGND sky130_fd_sc_hd__inv_2
X$12327 VGND \$1152 \$2329 \$1627 \$2306 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12328 VPWR VGND \$2049 \$294 \$2329 \$2306 \$2050 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12329 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12330 VPWR VGND \$2049 \$1179 \$2305 \$2272 \$2050 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12331 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12332 VGND \$1152 \$2305 \$2255 \$2272 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12334 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12335 VPWR VGND VPWR \$2287 \$1065 \$2330 \$1715 \$1955 VGND
+ sky130_fd_sc_hd__and4_1
X$12336 VPWR VGND VPWR \$2275 \$1914 \$1956 \$2219 \$2229 VGND
+ sky130_fd_sc_hd__and4_1
X$12337 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12338 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12339 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12340 VPWR VGND VPWR \$2146 \$2276 \$2287 \$2275 \$2273 VGND
+ sky130_fd_sc_hd__and4_1
X$12341 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12342 VPWR \$2348 VPWR VGND \$1128 \$1360 \$1705 VGND sky130_fd_sc_hd__or3_1
X$12343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12344 VGND \$2348 \$2357 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12345 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12346 VGND \$2288 \$2369 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12347 VPWR \$1448 \$2288 \$1415 VPWR VGND \$1360 \$1679 VGND
+ sky130_fd_sc_hd__or4_1
X$12348 VPWR \$2349 VPWR VGND \$1322 \$1449 \$1679 VGND sky130_fd_sc_hd__or3_1
X$12349 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12351 VGND \$2331 \$2330 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12352 VPWR \$2289 VGND \$2277 \$1782 VPWR VGND sky130_fd_sc_hd__or2_1
X$12353 VGND \$2289 \$2073 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12355 VGND \$2332 \$1957 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$12356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12357 VGND \$2241 \$1966 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12358 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12359 VGND \$358 \$2255 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12360 VGND \$2290 \$2043 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12362 VPWR VGND \$2401 \$1594 \$2333 \$2278 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12364 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12365 VPWR \$2324 \$2333 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12367 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12368 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12370 VPWR \$2307 \$2165 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12372 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12374 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12375 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12376 VGND \$1152 \$2350 \$2232 \$2308 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12377 VPWR VGND \$2127 \$354 \$2350 \$2308 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12380 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12383 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12384 VGND \$1152 \$2207 \$2232 \$2208 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12385 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12387 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12389 VPWR VGND \$2351 VPWR mgmt_gpio_in[6] VGND sky130_fd_sc_hd__buf_2
X$12390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12392 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12393 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12395 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12396 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12397 VPWR \$2422 \$2423 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12398 VPWR \$2387 VGND VPWR sram_ro_data[30] VGND sky130_fd_sc_hd__clkbuf_1
X$12399 VPWR \$2435 VGND \$2234 VPWR \$2194 VGND sky130_fd_sc_hd__nor2_1
X$12400 VPWR \$2388 VPWR VGND \$2424 \$1998 VGND sky130_fd_sc_hd__or2_2
X$12401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12403 VPWR \$2389 VGND \$2424 \$1963 VPWR VGND sky130_fd_sc_hd__or2_1
X$12404 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12405 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12406 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12407 VPWR VGND VPWR \$2352 \$2389 VGND sky130_fd_sc_hd__inv_2
X$12408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12409 VPWR \$2436 VGND \$2320 VPWR \$2194 VGND sky130_fd_sc_hd__nor2_1
X$12410 VPWR \$2623 \$2243 \$2436 VPWR VGND \$2409 \$2437 VGND
+ sky130_fd_sc_hd__or4_1
X$12411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12412 VPWR \$2437 VGND \$2234 VPWR \$1999 VGND sky130_fd_sc_hd__nor2_1
X$12413 VPWR \$2438 VGND \$2409 \$2468 VPWR VGND sky130_fd_sc_hd__or2_1
X$12414 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12416 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12417 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12418 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12419 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12420 VPWR \$2426 \$2411 \$2438 VPWR VGND \$2364 \$2425 VGND
+ sky130_fd_sc_hd__or4_1
X$12421 VPWR \$2469 \$2452 \$2353 VPWR VGND \$2354 \$2391 VGND
+ sky130_fd_sc_hd__or4_1
X$12422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12424 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12425 VPWR VGND \$2390 VPWR \$2412 \$2452 \$2439 VGND sky130_fd_sc_hd__a21o_1
X$12426 VPWR VGND \$2471 VPWR \$2412 \$2439 \$2470 VGND sky130_fd_sc_hd__a21o_1
X$12427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12428 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12429 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12430 VPWR VPWR \$2453 VGND \$2472 \$2427 \$1980 VGND sky130_fd_sc_hd__o21ai_1
X$12431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12432 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12433 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12434 VPWR \$2441 VPWR VGND \$2440 \$1887 \$2427 VGND sky130_fd_sc_hd__or3_1
X$12435 VPWR \$2428 VGND \$2440 \$2470 VPWR VGND sky130_fd_sc_hd__or2_1
X$12436 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12437 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12438 VPWR \$2442 VGND \$2392 \$2428 VPWR VGND sky130_fd_sc_hd__or2_1
X$12439 VGND \$2410 \$2444 \$2441 \$2413 \$2443 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$12440 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12441 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12442 VPWR \$2454 VGND \$2393 \$2442 VPWR VGND sky130_fd_sc_hd__or2_1
X$12443 VPWR \$2443 \$2427 VGND \$2411 VPWR \$2445 \$2414 VGND
+ sky130_fd_sc_hd__or4_2
X$12444 VPWR \$2489 VGND \$2394 \$2454 VPWR VGND sky130_fd_sc_hd__or2_1
X$12445 VPWR \$2682 VPWR VGND \$2553 \$2198 \$2414 VGND sky130_fd_sc_hd__or3_1
X$12446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12450 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12454 VGND \$856 \$2415 \$1750 \$2446 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12456 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12457 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12458 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12459 VPWR VGND \$2321 \$183 \$2415 \$2446 \$2322 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12460 VPWR \$2088 \$2415 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12465 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12466 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12467 VPWR VGND \$2120 \$281 \$2455 \$2491 \$2106 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12469 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12470 VPWR VGND \$2120 \$294 \$2473 \$2492 \$2106 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12473 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12474 VGND \$2429 \$1113 \$2524 \$2474 \$456 \$588 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12477 VPWR \$2475 VGND VPWR \$2323 \$1954 \$2342 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$12478 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12480 VPWR \$2476 VGND VPWR \$1325 \$2456 \$2072 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$12481 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12482 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12484 VGND \$2478 \$2476 \$1192 \$2525 \$2458 \$2477 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12488 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12489 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12490 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12492 VPWR VGND VPWR \$2459 \$2479 \$2478 \$2495 \$2371 VGND
+ sky130_fd_sc_hd__and4_1
X$12493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12495 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12496 VPWR \$1598 VGND VPWR \$2386 \$1454 VGND sky130_fd_sc_hd__or2_4
X$12497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12498 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12499 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12500 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12501 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12502 VPWR \$1598 VGND VPWR \$2497 \$1426 VGND sky130_fd_sc_hd__or2_4
X$12503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12504 VGND \$1947 \$2430 \$1645 \$1556 \$2422 \$2431 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$12505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12506 VPWR \$1598 VGND VPWR \$2375 \$1329 VGND sky130_fd_sc_hd__or2_4
X$12507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12508 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12511 VGND \$2499 \$762 \$2005 \$2500 \$2301 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$12512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12513 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12514 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12515 VGND \$2501 \$1792 \$2327 \$2065 \$2046 \$1240 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12519 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12520 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12522 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12523 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12525 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12526 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12527 VGND \$2504 \$2480 \$861 \$1953 \$1987 \$2324 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12530 VPWR \$2505 VGND VPWR \$1294 \$1793 \$1943 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$12531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12534 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12537 VPWR \$2461 VGND VPWR \$475 \$456 \$2481 \$2447 VGND
+ sky130_fd_sc_hd__o22a_1
X$12538 VGND \$1928 \$2395 \$2531 \$2375 \$2325 \$2432 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12539 VGND \$2482 \$2461 \$1702 \$1198 \$379 \$731 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12540 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12541 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12542 VPWR \$2448 VPWR VGND \$1128 \$1360 \$1679 VGND sky130_fd_sc_hd__or3_1
X$12543 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12545 VGND \$2448 \$2525 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12547 VGND \$2417 \$2458 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12549 VGND \$2418 \$2416 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12550 VPWR \$2508 VPWR VGND \$1384 \$1438 \$1705 VGND sky130_fd_sc_hd__or3_1
X$12551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12552 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12555 VPWR \$2462 VPWR VGND \$1438 \$1360 \$1705 VGND sky130_fd_sc_hd__or3_1
X$12556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12557 VPWR \$2519 VPWR VGND \$1322 \$1438 \$1705 VGND sky130_fd_sc_hd__or3_1
X$12558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12559 VPWR \$2463 VGND \$2325 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$12560 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12561 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12562 VGND \$2483 \$2590 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$12563 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12564 VPWR VGND \$2334 VPWR \$2463 VGND sky130_fd_sc_hd__clkbuf_4
X$12565 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12566 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12567 VPWR \$2432 \$2465 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12568 VPWR VGND \$2401 \$411 \$2465 \$2509 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12569 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12570 VGND \$1152 \$2465 \$2450 \$2509 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12571 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12572 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12573 VPWR VGND \$2401 \$542 \$2402 \$2419 \$2334 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12574 VGND \$1152 \$2402 \$2450 \$2419 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12576 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12577 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12578 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12579 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12580 VGND \$1152 \$2404 \$2232 \$2420 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12581 VPWR VGND VPWR \$2464 \$2404 VGND sky130_fd_sc_hd__inv_2
X$12582 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12583 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12584 VGND \$1152 \$2466 \$2232 \$2484 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12585 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12586 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12587 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12588 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12589 VPWR VGND VPWR \$2449 \$2379 VGND sky130_fd_sc_hd__inv_2
X$12590 VPWR VGND \$2127 \$1594 \$2433 \$2451 \$2128 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12591 VPWR \$2460 \$2433 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12592 VGND \$1152 \$2433 \$2232 \$2451 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12593 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12594 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12595 VPWR \$2405 VGND VPWR \$2403 VGND sky130_fd_sc_hd__clkbuf_1
X$12596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12597 VPWR VGND mgmt_gpio_oeb[6] VPWR \$2421 VGND sky130_fd_sc_hd__buf_2
X$12598 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12604 VGND spi_csb \$3321 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$12605 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12606 VPWR \$3300 VPWR VGND \$2320 VGND sky130_fd_sc_hd__buf_4
X$12607 VPWR \$3300 VGND \$2015 \$3342 VPWR VGND sky130_fd_sc_hd__or2_1
X$12608 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12609 VPWR VPWR \$3322 VGND \$2996 \$1998 \$2336 \$3057 VGND
+ sky130_fd_sc_hd__a211o_1
X$12610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12611 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12613 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12614 VPWR VGND \$3341 VPWR \$3359 \$3358 \$3340 VGND sky130_fd_sc_hd__a21o_1
X$12615 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12616 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12618 VPWR VGND \$1999 VPWR \$3299 VGND sky130_fd_sc_hd__clkbuf_4
X$12619 VGND \$3256 \$2640 \$2001 \$2537 \$3341 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2bb2o_1
X$12620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12621 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12622 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12623 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12624 VPWR VGND VPWR \$3301 \$3258 VGND sky130_fd_sc_hd__inv_2
X$12625 VGND \$2942 \$2891 \$2931 \$3638 \$3301 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$12626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12628 VPWR VGND \$2891 VPWR \$3360 VGND sky130_fd_sc_hd__clkbuf_4
X$12629 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12630 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12632 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12636 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12637 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12638 VPWR \$3361 VGND \$3141 VPWR \$3342 VGND sky130_fd_sc_hd__nor2_1
X$12639 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12640 VGND \$3302 \$3323 \$3261 \$2950 \$2445 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$12641 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12642 VPWR \$3443 VGND \$3361 \$3179 VPWR VGND sky130_fd_sc_hd__or2_1
X$12643 VPWR \$3261 VPWR VGND \$2663 \$3343 \$3361 VGND sky130_fd_sc_hd__or3_2
X$12644 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12645 VPWR \$3362 VGND \$3282 \$3343 VPWR VGND sky130_fd_sc_hd__or2_1
X$12646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12647 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12649 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12650 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12651 VGND \$2777 \$3305 \$2556 \$3303 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12652 VPWR VPWR VGND \$3324 \$3126 VGND sky130_fd_sc_hd__clkbuf_2
X$12653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12654 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12655 VPWR VGND \$3284 \$293 \$3305 \$3303 \$3304 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12656 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12657 VPWR VGND \$3284 \$294 \$3270 \$3283 \$3304 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12658 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12659 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12660 VGND \$856 \$3285 \$2556 \$3306 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12661 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12662 VPWR VPWR VGND \$3344 \$3304 VGND sky130_fd_sc_hd__clkbuf_2
X$12663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12664 VPWR \$3344 VGND \$2314 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$12665 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12667 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12668 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12669 VPWR VPWR VGND \$3286 \$3324 VGND sky130_fd_sc_hd__clkbuf_2
X$12670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12671 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12672 VPWR VPWR VGND \$3133 \$3363 VGND sky130_fd_sc_hd__clkbuf_2
X$12673 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12675 VPWR VGND VPWR \$3217 \$3345 VGND sky130_fd_sc_hd__inv_2
X$12676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12678 VPWR \$1435 VGND VPWR \$3042 \$1571 VGND sky130_fd_sc_hd__or2_4
X$12679 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12680 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12681 VGND \$3308 \$3346 \$2609 \$2330 \$2219 \$3333 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12682 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12683 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12684 VPWR \$1103 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12685 VGND \$3365 \$3347 \$1017 \$1103 \$1219 \$3364 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12687 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12688 VGND \$3309 \$2218 \$3348 \$1065 \$880 \$3132 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12689 VPWR \$2099 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12690 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12692 VGND \$3310 \$2227 \$868 \$2073 \$2096 \$3349 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12693 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12694 VPWR \$2099 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12695 VPWR VGND VPWR \$3325 \$3310 \$3308 \$3309 \$2099 VGND
+ sky130_fd_sc_hd__and4_1
X$12696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12697 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12698 VPWR \$488 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12699 VPWR \$3334 VGND VPWR \$3333 \$3042 \$488 \$326 VGND
+ sky130_fd_sc_hd__o22a_1
X$12700 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12701 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12702 VGND \$3366 \$3334 \$712 \$1266 \$1466 \$3417 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12703 VGND \$3311 \$725 \$1266 \$1219 \$3312 \$1657 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$12704 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12706 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12707 VGND \$3289 \$3367 \$2060 \$2355 \$1819 \$3350 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12708 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12709 VPWR \$3326 VGND VPWR \$3180 \$2372 \$3265 \$2497 VGND
+ sky130_fd_sc_hd__o22a_1
X$12710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12712 VPWR \$881 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12713 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12714 VGND \$3288 \$881 \$3351 \$2386 \$2314 \$3508 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12715 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12716 VGND mgmt_gpio_in[4] \$3286 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12718 VGND \$3370 \$3326 \$3368 \$2614 \$1300 \$1617 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12719 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12720 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12722 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12723 VPWR \$2114 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12724 VGND \$3371 \$3369 \$424 \$1953 \$1987 \$3263 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12726 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12727 VPWR \$2114 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$12728 VPWR VGND VPWR \$3335 \$3373 \$3206 \$3372 \$2181 VGND
+ sky130_fd_sc_hd__and4_1
X$12729 VPWR VGND VPWR \$3327 \$2114 \$3314 \$3291 \$3313 VGND
+ sky130_fd_sc_hd__and4_1
X$12730 VPWR \$3696 VGND VPWR \$424 \$2045 \$3061 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$12731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12733 VPWR \$3374 VGND VPWR \$3352 \$2919 \$1602 \$1890 VGND
+ sky130_fd_sc_hd__o22a_1
X$12734 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12735 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12736 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12739 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12740 VPWR \$3376 VGND VPWR \$576 \$2045 \$2994 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$12741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12742 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12743 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12744 VGND \$3377 \$3330 \$576 \$1953 \$1987 \$2360 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12745 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12748 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12749 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12750 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12752 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12754 VGND \$3293 \$3315 \$731 \$1953 \$1987 \$2432 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12755 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12757 VGND \$4109 \$3316 \$3274 \$3064 VPWR \$821 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$12758 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12759 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12760 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12761 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12762 VPWR \$3379 VGND VPWR \$1720 \$1776 \$1557 \$1743 VGND
+ sky130_fd_sc_hd__o22a_1
X$12763 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12764 VGND \$3337 \$3353 \$385 \$1953 \$1987 \$3294 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12766 VPWR \$3380 VGND VPWR \$385 \$2045 \$2976 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$12767 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12768 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12770 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12771 VGND \$3381 \$3354 \$2005 \$3355 \$3337 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$12772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12774 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12775 VPWR \$3382 VGND VPWR \$2053 \$2180 \$3338 \$1839 VGND
+ sky130_fd_sc_hd__o22a_1
X$12776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12777 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12778 VGND \$3383 \$3382 \$3354 \$1879 \$2785 \$2976 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$12779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12781 VPWR \$3351 \$3317 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12782 VPWR VGND \$2633 \$386 \$3317 \$3318 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12783 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12784 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12785 VGND \$2989 \$3317 \$2450 \$3318 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12786 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12789 VPWR VGND \$2694 \$1179 \$3385 \$3386 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12790 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12792 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12793 VGND \$2989 \$3296 \$2232 \$3295 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12794 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12795 VPWR VGND VPWR \$3338 \$3296 VGND sky130_fd_sc_hd__inv_2
X$12796 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12798 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12799 VPWR VGND \$3319 \$2829 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$12800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12801 VPWR VGND \$3169 \$184 \$3331 \$3320 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12802 VGND \$1152 \$3331 \$2232 \$3320 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12803 VPWR \$3242 \$3331 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12804 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12805 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12806 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12807 VPWR \$3387 VGND VPWR mgmt_gpio_in[9] VGND sky130_fd_sc_hd__clkbuf_1
X$12808 VPWR VGND VPWR \$3352 \$3387 VGND sky130_fd_sc_hd__inv_2
X$12809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12810 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12811 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12814 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12815 VGND \$4601 \$4651 \$4879 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$12816 VPWR VGND wb_dat_o[19] VPWR \$4907 VGND sky130_fd_sc_hd__buf_2
X$12817 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12819 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12820 VPWR \$4833 \$4842 \$4881 VPWR VGND \$4891 \$4880 VGND
+ sky130_fd_sc_hd__or4_1
X$12821 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12822 VGND \$4880 \$2537 \$4891 \$4881 \$4864 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$12823 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12824 VPWR \$4833 VPWR VGND \$3916 \$4891 \$4880 VGND sky130_fd_sc_hd__or3_2
X$12825 VPWR \$4908 VPWR VGND \$3057 VGND sky130_fd_sc_hd__buf_4
X$12826 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12827 VGND \$4881 \$3299 \$4833 \$4853 \$4863 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$12828 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12829 VGND \$3410 \$4916 \$4941 \$4687 \$4909 \$4075 VPWR VPWR VGND
+ sky130_fd_sc_hd__a41o_2
X$12830 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12831 VPWR VPWR VGND \$4266 \$4651 VGND sky130_fd_sc_hd__clkbuf_2
X$12832 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12834 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12835 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12836 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12837 VGND \$4853 \$2337 \$4863 \$4881 \$4864 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$12838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12839 VPWR \$4891 \$4902 \$4853 VPWR VGND \$4833 \$4881 VGND
+ sky130_fd_sc_hd__or4_1
X$12840 VPWR \$4249 VPWR VGND \$4892 \$4833 VGND sky130_fd_sc_hd__or2_2
X$12841 VPWR VGND VPWR \$4577 \$4910 VGND sky130_fd_sc_hd__inv_2
X$12842 VPWR VPWR \$4917 VGND \$4910 \$4919 \$3919 VGND sky130_fd_sc_hd__o21ai_1
X$12843 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12844 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12845 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12846 VGND \$4663 \$4918 \$3857 \$4664 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$12847 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12848 VPWR VGND VPWR \$4931 \$3155 VGND sky130_fd_sc_hd__inv_2
X$12849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12850 VGND \$4920 \$4931 \$4597 \$4664 \$4911 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$12851 VPWR \$4911 VGND \$4919 \$4578 VPWR VGND sky130_fd_sc_hd__or2_1
X$12852 VPWR \$4663 VPWR \$4597 \$4903 VGND \$4326 \$4893 \$4664 VGND
+ sky130_fd_sc_hd__a311oi_1
X$12853 VPWR \$4894 VGND \$4920 \$4855 VPWR VGND sky130_fd_sc_hd__or2_1
X$12854 VPWR \$4893 VGND \$4894 \$4800 VPWR VGND sky130_fd_sc_hd__or2_1
X$12855 VPWR \$4664 \$4603 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12856 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12857 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12858 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12860 VPWR VPWR \$4181 VGND \$4912 \$2640 \$4736 \$4882 VGND
+ sky130_fd_sc_hd__a211o_1
X$12861 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12863 VPWR \$4819 VGND \$4895 VPWR \$3892 VGND sky130_fd_sc_hd__nor2_1
X$12864 VPWR \$4883 VGND \$4895 VPWR \$2996 VGND sky130_fd_sc_hd__nor2_1
X$12865 VGND \$1963 \$4895 \$1998 \$4895 \$4553 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22ai_4
X$12866 VPWR \$4866 VGND \$4883 \$4153 VPWR VGND sky130_fd_sc_hd__or2_1
X$12867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12868 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12870 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12872 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12874 VPWR \$4904 VGND \$4932 \$4820 VPWR VGND sky130_fd_sc_hd__or2_1
X$12875 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12876 VPWR \$4886 VPWR VGND \$4896 \$4868 VGND sky130_fd_sc_hd__nand2_1
X$12877 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12879 VPWR \$4904 VGND \$4913 VPWR \$4869 VGND sky130_fd_sc_hd__or2b_1
X$12880 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12881 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12884 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12886 VGND \$3272 \$4897 \$4159 \$1369 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$12887 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12888 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12889 VPWR VGND \$4701 \$3732 \$4923 \$4922 \$4677 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12890 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12892 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12893 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12894 VPWR VGND VPWR \$2819 \$4923 VGND sky130_fd_sc_hd__inv_2
X$12895 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12897 VPWR VGND \$4760 \$3711 \$4845 \$4870 \$4717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12898 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12900 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12901 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12907 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12908 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12910 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12911 VPWR \$4654 \$4667 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12912 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12914 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12915 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12916 VGND \$4761 \$4847 \$4813 \$4898 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12918 VPWR VGND \$4899 \$4023 \$4847 \$4898 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12920 VPWR VGND \$4899 \$3711 \$4848 \$4872 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12921 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12922 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12927 VPWR VGND \$4899 \$1179 \$4874 \$4873 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12928 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12929 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12930 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12931 VGND \$4353 \$4824 \$4850 \$4887 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12932 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12933 VPWR VGND \$4899 \$1594 \$4824 \$4887 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12935 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12936 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12937 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12938 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12940 VPWR VGND \$4905 \$1594 \$4901 \$4914 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12941 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12942 VPWR VGND VPWR \$2286 \$4901 VGND sky130_fd_sc_hd__inv_2
X$12943 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12944 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12945 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12946 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12947 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12950 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12953 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12954 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12955 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12956 VGND \$3952 \$4765 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$12957 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12958 VGND \$4764 \$4876 \$4765 \$4888 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$12959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12960 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12961 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12963 VPWR VGND \$4905 \$184 \$4925 \$4924 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12964 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12965 VPWR VGND \$5100 VPWR \$4889 VGND sky130_fd_sc_hd__clkbuf_4
X$12966 VPWR \$3678 \$4925 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$12967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12969 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12971 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12972 VGND \$4353 \$4851 \$4427 \$4915 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$12973 VPWR VGND \$4709 \$1171 \$4851 \$4915 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12976 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$12977 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12978 VPWR VGND \$4709 \$3694 \$4877 \$4906 \$4710 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$12979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12980 VGND \$4353 \$4877 \$4828 \$4906 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$12981 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12982 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12983 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12984 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12986 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$12989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12990 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12992 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12993 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12994 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$12995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$12996 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$12997 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$12998 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$12999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13000 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13001 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13002 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13003 VPWR VGND wb_dat_o[27] VPWR \$5243 VGND sky130_fd_sc_hd__buf_2
X$13004 VGND \$4949 \$4651 \$5256 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$13005 VGND \$5256 \$4949 \$5076 \$5077 \$2221 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$13006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13008 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13009 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13010 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13011 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13012 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13013 VPWR \$4193 VPWR VGND \$5268 \$4474 VGND sky130_fd_sc_hd__or2_2
X$13014 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13016 VPWR \$5244 VGND \$3892 \$5147 VPWR VGND sky130_fd_sc_hd__or2_1
X$13017 VGND \$5244 \$2552 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$13018 VPWR VGND VPWR \$4818 \$5268 VGND sky130_fd_sc_hd__inv_2
X$13019 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13020 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13022 VPWR \$5190 VPWR VGND \$4833 \$4733 \$5274 VGND sky130_fd_sc_hd__or3_1
X$13023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13024 VPWR VPWR VGND \$4854 \$5245 \$4733 \$5274 VGND sky130_fd_sc_hd__a21o_2
X$13025 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13026 VPWR \$5170 VGND \$5245 VPWR \$4864 VGND sky130_fd_sc_hd__nor2_1
X$13027 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13029 VPWR \$5040 VPWR VGND \$5274 \$4930 \$4917 VGND sky130_fd_sc_hd__or3_2
X$13030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13031 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13032 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13033 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13034 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13035 VPWR \$4818 VPWR \$5269 VGND \$5220 \$4615 VGND sky130_fd_sc_hd__o21a_1
X$13036 VPWR \$5257 VGND \$2552 \$4698 VPWR VGND sky130_fd_sc_hd__or2_1
X$13037 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13039 VPWR VGND VPWR \$4615 \$5257 VGND sky130_fd_sc_hd__inv_2
X$13040 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13041 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13042 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13043 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13046 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13047 VPWR VGND VPWR \$5259 \$5290 VGND sky130_fd_sc_hd__inv_2
X$13048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13049 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13050 VGND \$4522 \$5258 \$5213 \$5259 \$5234 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$13051 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13052 VPWR \$5275 VPWR VGND \$5183 \$5269 \$5223 VGND sky130_fd_sc_hd__or3_1
X$13053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13055 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13057 VPWR \$5202 VPWR VGND \$4676 \$4727 \$5246 VGND sky130_fd_sc_hd__or3_1
X$13058 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13059 VPWR VGND \$5247 \$5246 \$4727 VPWR \$4582 \$5286 VGND
+ sky130_fd_sc_hd__or4b_2
X$13060 VPWR \$5223 VGND \$5247 \$4758 VPWR VGND sky130_fd_sc_hd__or2_1
X$13061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13062 VPWR \$4896 VGND \$5276 \$5246 VPWR VGND sky130_fd_sc_hd__or2_1
X$13063 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13064 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13065 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13067 VPWR \$5248 VGND VPWR \$5236 VGND sky130_fd_sc_hd__clkbuf_1
X$13068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13069 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13071 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13072 VPWR \$5260 VGND \$5184 VPWR \$5270 VGND sky130_fd_sc_hd__nor2_1
X$13073 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13074 VPWR VPWR VGND \$4715 \$5034 VGND sky130_fd_sc_hd__clkbuf_2
X$13075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13076 VPWR VGND VPWR \$5224 \$5226 VGND sky130_fd_sc_hd__inv_2
X$13077 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13079 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13080 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13081 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13082 VGND \$2777 \$5227 \$5165 \$5249 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13084 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13085 VPWR VGND \$5118 \$4774 \$5227 \$5249 \$5080 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13087 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13088 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13089 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13090 VGND \$4761 \$5228 \$5165 \$5237 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$13091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13092 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13093 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13094 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13096 VPWR VGND \$5097 \$411 \$5277 \$5287 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13099 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13100 VGND \$4774 \$1179 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$13101 VPWR VGND VPWR \$3842 \$5250 VGND sky130_fd_sc_hd__inv_2
X$13102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13103 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13105 VPWR VGND \$5229 \$1594 \$5193 \$5206 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13108 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13109 VGND \$4761 \$5217 \$4994 \$5216 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13113 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13114 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13115 VGND \$4761 \$5230 \$4994 \$5261 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13117 VPWR VGND \$5252 \$1594 \$5230 \$5261 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13118 VPWR VGND \$5262 VPWR \$5240 VGND sky130_fd_sc_hd__clkbuf_4
X$13119 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13121 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13122 VGND \$4761 \$5231 \$4850 \$5241 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13123 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13124 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13126 VPWR VGND \$5252 \$386 \$5194 \$5208 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13131 VGND \$4761 \$5253 \$4850 \$5271 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13133 VPWR VGND \$5252 \$411 \$5253 \$5271 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13135 VPWR \$5263 VGND \$1845 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$13136 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13137 VPWR VGND VPWR \$4319 \$5253 VGND sky130_fd_sc_hd__inv_2
X$13138 VPWR \$4123 \$5277 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13139 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13140 VGND \$4761 \$5254 \$5272 \$5273 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13141 VPWR VGND \$5044 \$411 \$5254 \$5273 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13142 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13143 VPWR \$5264 VGND \$2447 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$13144 VPWR VGND \$5086 \$184 \$5255 \$5242 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13145 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13146 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13148 VGND \$4764 \$5255 \$5006 \$5242 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13149 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13150 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13152 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13154 VPWR VGND VPWR \$5044 \$5035 VGND sky130_fd_sc_hd__inv_2
X$13155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13157 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13159 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13160 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13161 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13162 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13163 VPWR \$5265 VGND \$4239 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$13164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13167 VPWR VGND \$5046 \$1171 \$5198 \$5232 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13170 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13174 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13175 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13176 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13177 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13179 VPWR VGND \$5266 VPWR \$4749 VGND sky130_fd_sc_hd__clkbuf_4
X$13180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13183 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13184 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13190 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13191 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13192 VPWR \$5278 VGND VPWR \$2866 VGND sky130_fd_sc_hd__clkbuf_1
X$13193 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13194 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13196 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13199 VPWR VGND wb_dat_o[30] VPWR \$5358 VGND sky130_fd_sc_hd__buf_2
X$13200 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13201 VPWR \$5374 VGND VPWR \$5024 \$5076 \$1769 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$13202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13204 VPWR \$5316 VGND VPWR \$5059 \$5076 \$1619 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$13205 VPWR \$5076 \$5077 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13206 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13207 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13208 VGND \$5059 \$4651 \$5316 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$13209 VPWR VGND \$5077 VPWR \$5360 VGND sky130_fd_sc_hd__clkbuf_4
X$13210 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13211 VPWR VGND VPWR \$4917 \$4942 VGND sky130_fd_sc_hd__inv_2
X$13212 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13213 VPWR \$4806 VGND \$5268 VPWR \$5326 VGND sky130_fd_sc_hd__nor2_1
X$13214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13215 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13216 VPWR \$5281 \$5386 \$4916 VPWR VGND \$4930 \$4917 VGND
+ sky130_fd_sc_hd__or4_1
X$13217 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13218 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13220 VPWR \$5375 VPWR VGND \$5025 \$4917 \$5359 VGND sky130_fd_sc_hd__or3_1
X$13221 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13222 VGND \$5219 \$5220 \$5285 \$5359 \$4930 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4b_1
X$13223 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13225 VGND \$5348 \$2471 \$5220 \$5457 \$4918 \$5361 VPWR VPWR VGND
+ sky130_fd_sc_hd__a311o_1
X$13226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13227 VPWR VPWR \$5257 VGND \$5326 \$5349 \$4807 VGND sky130_fd_sc_hd__o21ai_1
X$13228 VPWR \$5221 VGND \$4918 \$5376 VPWR VGND sky130_fd_sc_hd__or2_1
X$13229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13231 VPWR \$5327 VGND \$5349 \$5350 VPWR VGND sky130_fd_sc_hd__or2_1
X$13232 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13233 VPWR \$5336 VGND \$5327 \$5328 VPWR VGND sky130_fd_sc_hd__or2_1
X$13234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13236 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13237 VPWR \$2683 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13239 VPWR \$2683 \$5293 \$5327 VPWR VGND \$5348 \$5290 VGND
+ sky130_fd_sc_hd__or4_1
X$13240 VPWR \$3323 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13242 VPWR \$3323 \$5362 \$5350 VPWR VGND \$5440 \$5328 VGND
+ sky130_fd_sc_hd__or4_1
X$13243 VPWR \$5362 \$5377 \$5361 VPWR VGND \$5304 \$5282 VGND
+ sky130_fd_sc_hd__or4_1
X$13244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13246 VPWR \$5337 VGND \$5377 \$5285 VPWR VGND sky130_fd_sc_hd__or2_1
X$13247 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13249 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13251 VPWR \$5294 VGND \$5337 \$4520 VPWR VGND sky130_fd_sc_hd__or2_1
X$13252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13253 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13254 VPWR \$5360 VGND \$5351 \$5235 VPWR VGND sky130_fd_sc_hd__or2_1
X$13255 VPWR \$5363 VGND \$5317 \$5235 VPWR VGND sky130_fd_sc_hd__or2_1
X$13256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13257 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13259 VPWR \$5329 VGND \$5305 \$5115 VPWR VGND sky130_fd_sc_hd__or2_1
X$13260 VGND \$5338 \$5329 \$3831 \$5318 \$4933 \$5301 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$13261 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13263 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13264 VPWR \$5306 VGND \$5184 VPWR \$5339 VGND sky130_fd_sc_hd__nor2_1
X$13265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13266 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13268 VPWR VPWR \$5339 VGND \$1315 \$5378 \$5351 VGND sky130_fd_sc_hd__o21ai_1
X$13269 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13270 VPWR VGND VPWR \$5351 \$5215 VGND sky130_fd_sc_hd__inv_2
X$13271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13272 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13273 VGND \$2777 \$5307 \$4811 \$5340 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13274 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13276 VPWR VGND \$5192 \$3711 \$5307 \$5340 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13278 VPWR VGND \$5118 \$3711 \$5341 \$5379 \$5080 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13280 VPWR VGND \$5118 \$4023 \$5330 \$5352 \$5080 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13281 VGND \$4761 \$5330 \$5165 \$5352 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13282 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13283 VGND \$3711 \$386 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$13284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13286 VPWR VGND VPWR \$3704 \$5330 VGND sky130_fd_sc_hd__inv_2
X$13287 VPWR VGND \$5097 \$354 \$5380 \$5381 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13288 VPWR VGND VPWR \$3961 \$5341 VGND sky130_fd_sc_hd__inv_2
X$13289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13290 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13291 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13292 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13293 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13294 VPWR VGND \$5380 \$3782 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13297 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13298 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13299 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13300 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13301 VPWR VGND \$5229 \$1171 \$5364 \$5382 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13302 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13303 VPWR VGND \$5229 \$386 \$5308 \$5342 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13305 VGND \$4761 \$5308 \$4994 \$5342 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13306 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13307 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13309 VPWR VGND \$5365 \$2804 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13310 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13311 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13312 VPWR VGND VPWR \$4544 \$5331 VGND sky130_fd_sc_hd__inv_2
X$13313 VGND \$4761 \$5343 \$4994 \$5353 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13315 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13316 VPWR VGND \$5252 \$4774 \$5343 \$5353 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13317 VGND \$4761 \$5331 \$5367 \$5366 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13318 VPWR VGND VPWR \$3399 \$5343 VGND sky130_fd_sc_hd__inv_2
X$13319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13321 VPWR VGND VPWR \$2647 \$5319 VGND sky130_fd_sc_hd__inv_2
X$13322 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13323 VPWR VGND \$5332 \$1594 \$5319 \$5354 \$5391 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13324 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13325 VGND \$4761 \$5319 \$5367 \$5354 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13328 VPWR VGND VPWR \$3673 \$5368 VGND sky130_fd_sc_hd__inv_2
X$13329 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13330 VGND \$4761 \$5309 \$5369 \$5370 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13331 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13332 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13333 VPWR VGND \$5252 \$354 \$5309 \$5370 \$5262 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13335 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13337 VGND \$4761 \$5310 \$5272 \$5320 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13338 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13339 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13341 VGND \$4761 \$5333 \$5272 \$5383 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13342 VPWR VGND \$5391 VPWR \$4693 VGND sky130_fd_sc_hd__clkbuf_4
X$13343 VPWR VGND VPWR \$4627 \$5333 VGND sky130_fd_sc_hd__inv_2
X$13344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13345 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13347 VPWR VGND \$5371 \$3476 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13348 VGND \$4764 \$5311 \$5334 \$5321 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13350 VPWR VGND VPWR \$3480 \$5372 VGND sky130_fd_sc_hd__inv_2
X$13351 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13352 VPWR VGND \$5344 \$354 \$5313 \$5322 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13353 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13355 VGND \$4764 \$5313 \$5334 \$5322 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13357 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13358 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13359 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13361 VPWR VGND \$5345 \$4774 \$5297 \$5314 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13365 VGND \$5296 \$4562 mgmt_gpio_out[33] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$13366 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13367 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13369 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13370 VPWR VGND \$5335 \$354 \$5299 \$5288 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13371 VPWR VGND VPWR \$5373 \$4724 VGND sky130_fd_sc_hd__inv_2
X$13372 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13373 VPWR VGND \$5335 \$1171 \$5324 \$5315 \$5266 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13375 VPWR VGND VPWR \$5335 \$5266 VGND sky130_fd_sc_hd__inv_2
X$13376 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13379 VGND \$5355 \$1171 \$5324 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13380 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13381 VPWR \$5356 VGND VPWR \$5355 \$4724 \$5325 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$13382 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13383 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13384 VGND \$5325 \$2866 mgmt_gpio_out[16] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$13385 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13386 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13389 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13390 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13393 VPWR \$2153 VGND VPWR sram_ro_data[27] VGND sky130_fd_sc_hd__clkbuf_1
X$13394 VPWR \$2210 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$13395 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13396 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13397 VPWR \$2154 VPWR VGND \$2015 \$2194 VGND sky130_fd_sc_hd__or2_2
X$13398 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13399 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13400 VPWR \$2195 VGND \$2154 \$1998 VPWR VGND sky130_fd_sc_hd__or2_1
X$13401 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13404 VPWR \$2213 VGND \$2212 \$2233 VPWR \$2222 VGND sky130_fd_sc_hd__and3b_1
X$13405 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13406 VPWR \$2234 VPWR \$2155 VGND \$2168 \$1999 VGND sky130_fd_sc_hd__o21a_1
X$13407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13409 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13410 VPWR VGND VPWR \$2235 \$2130 VGND sky130_fd_sc_hd__inv_2
X$13411 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13413 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13414 VPWR \$2236 VPWR VGND \$2243 \$2235 \$2311 VGND sky130_fd_sc_hd__or3_1
X$13415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13416 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13417 VPWR \$1899 VGND \$2234 VPWR \$2002 VGND sky130_fd_sc_hd__nor2_1
X$13418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13420 VGND \$2215 \$2213 \$2196 \$2223 \$1977 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4b_4
X$13421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13423 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13424 VPWR VGND \$1897 \$2257 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13426 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13427 VGND \$2216 \$2171 \$2224 \$2214 \$2027 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$13428 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13429 VGND \$2189 \$2257 \$2171 \$2214 \$2058 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$13430 VPWR \$2258 VGND \$2237 \$2259 VPWR VGND sky130_fd_sc_hd__or2_1
X$13431 VPWR \$2259 VGND \$2026 VPWR \$1963 VGND sky130_fd_sc_hd__nor2_1
X$13432 VPWR \$2237 VGND \$2216 \$2104 VPWR VGND sky130_fd_sc_hd__or2_1
X$13433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13434 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13435 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13436 VPWR \$2238 VGND \$2173 \$2217 VPWR VGND sky130_fd_sc_hd__or2_1
X$13437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13439 VPWR VGND \$1725 \$2244 \$2261 \$2260 \$1712 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13442 VGND \$856 \$2199 \$1750 \$2245 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13444 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13445 VGND \$463 \$1750 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$13446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13448 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13450 VGND \$463 \$3030 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$13451 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13456 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13458 VPWR VGND VPWR \$2225 \$2158 VGND sky130_fd_sc_hd__inv_2
X$13459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13461 VPWR VGND \$2120 \$293 \$2263 \$2262 \$2106 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13464 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13465 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13466 VPWR \$2246 VGND \$2190 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$13467 VPWR VPWR VGND \$2246 \$2106 VGND sky130_fd_sc_hd__clkbuf_2
X$13468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13470 VPWR \$2264 VGND VPWR \$1163 \$2135 \$1744 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$13471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13473 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13474 VPWR VGND VPWR \$2268 \$2267 \$2265 \$2266 \$2228 VGND
+ sky130_fd_sc_hd__and4_1
X$13475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13477 VGND \$2248 \$2268 \$2269 VPWR \$526 VPWR VGND sky130_fd_sc_hd__nand3_4
X$13478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13480 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13481 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13484 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13486 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13487 VPWR \$2239 VGND VPWR \$1744 \$1967 \$2225 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$13488 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13489 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13491 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13492 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13494 VPWR \$2270 VGND VPWR \$2292 \$1967 \$2176 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$13495 VPWR \$2271 VGND VPWR \$920 \$1421 \$2176 \$1713 VGND
+ sky130_fd_sc_hd__o22a_1
X$13496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13497 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13498 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13499 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13500 VGND \$2249 \$1024 \$1421 \$2180 \$2191 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$13501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13503 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13504 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13506 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13508 VPWR \$2250 VGND VPWR \$920 \$1956 \$1778 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$13509 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13511 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13512 VPWR \$2251 VGND VPWR \$1284 \$1421 \$2252 \$1867 VGND
+ sky130_fd_sc_hd__o22a_1
X$13513 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13516 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13518 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13519 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13520 VPWR \$464 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13521 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13522 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13523 VPWR \$2253 VGND \$2113 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$13524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13525 VPWR VPWR VGND \$2253 \$2050 VGND sky130_fd_sc_hd__clkbuf_2
X$13526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13528 VPWR VGND VPWR \$2273 \$2096 \$1966 \$2048 \$2007 VGND
+ sky130_fd_sc_hd__and4_1
X$13529 VPWR VGND VPWR \$2276 \$2358 \$2274 \$2254 \$2047 VGND
+ sky130_fd_sc_hd__and4_1
X$13530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13531 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13534 VGND \$2201 \$2226 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13536 VGND \$2183 \$2219 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13537 VGND \$2230 \$2274 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13538 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13539 VGND \$2240 \$2229 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13540 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13541 VPWR \$2240 VPWR VGND \$1814 \$1663 \$1782 VGND sky130_fd_sc_hd__or3_1
X$13542 VPWR \$2230 VPWR VGND \$1814 \$1797 \$1782 VGND sky130_fd_sc_hd__or3_1
X$13543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13544 VPWR \$2277 VGND \$1783 \$1797 VPWR VGND sky130_fd_sc_hd__or2_1
X$13545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13546 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13547 VPWR \$2241 VGND \$2231 \$1780 VPWR VGND sky130_fd_sc_hd__or2_1
X$13548 VPWR \$2231 VGND \$1783 \$1663 VPWR VGND sky130_fd_sc_hd__or2_1
X$13549 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13550 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13551 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13552 VPWR \$2242 VGND \$1782 \$1531 VPWR VGND sky130_fd_sc_hd__or2_1
X$13553 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13554 VGND \$2242 \$2254 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13555 VGND \$2202 \$2107 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13556 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13558 VGND \$1152 \$2333 \$2255 \$2278 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13559 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13560 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13561 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13562 VPWR VGND VPWR \$2191 \$2203 VGND sky130_fd_sc_hd__inv_2
X$13563 VGND \$1152 \$2203 \$1273 \$2204 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13565 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13566 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13567 VGND \$1152 \$2165 \$2232 \$2150 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13568 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13569 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13572 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13573 VPWR VGND VPWR \$2252 \$2205 VGND sky130_fd_sc_hd__inv_2
X$13574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13576 VGND \$1152 \$2205 \$2232 \$2206 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13577 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13578 VPWR VGND VPWR \$2127 \$2128 VGND sky130_fd_sc_hd__inv_2
X$13579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13580 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13581 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13582 VPWR VGND \$2207 \$2033 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13583 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13584 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13586 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13587 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13590 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13592 VPWR \$1496 \$1112 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13594 VPWR \$1451 \$1459 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13595 VGND \$1499 \$1498 \$381 \$1497 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$13596 VPWR \$1459 VGND VPWR sram_ro_data[15] VGND sky130_fd_sc_hd__clkbuf_1
X$13597 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13598 VPWR \$1472 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$13599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13600 VPWR \$1499 VGND VPWR \$1472 VGND sky130_fd_sc_hd__clkbuf_1
X$13601 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13604 VPWR VGND \$1473 VPWR \$1279 VGND sky130_fd_sc_hd__clkbuf_4
X$13605 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13607 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13608 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13613 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13614 VPWR \$1500 VPWR VGND \$1433 \$1485 VGND sky130_fd_sc_hd__nand2_1
X$13615 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13616 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13617 VGND \$1442 \$1487 \$1461 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13618 VPWR \$1485 VPWR \$1461 VGND \$1500 \$1433 VGND sky130_fd_sc_hd__o21a_1
X$13619 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13620 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13621 VPWR VGND VPWR \$1485 \$1486 VGND sky130_fd_sc_hd__inv_2
X$13622 VPWR \$1386 VPWR \$1501 VGND \$1486 \$1487 VGND sky130_fd_sc_hd__o21a_1
X$13623 VPWR \$1486 VPWR VGND \$1487 \$1386 VGND sky130_fd_sc_hd__nand2_1
X$13624 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13626 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13627 VGND \$1502 \$1337 \$1487 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13629 VGND \$1462 \$1502 \$1488 \$1369 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$13630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13631 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13632 VPWR VGND \$1525 VPWR \$1504 \$1503 \$1453 VGND sky130_fd_sc_hd__a21o_1
X$13633 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13635 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13636 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13639 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13641 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13642 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13646 VPWR \$1463 VPWR VGND \$1489 \$1474 \$1526 VGND sky130_fd_sc_hd__or3_1
X$13647 VPWR \$1475 VPWR VGND \$1462 \$1474 \$1453 VGND sky130_fd_sc_hd__or3_1
X$13648 VPWR \$1476 VPWR VGND \$1489 \$1474 \$1453 VGND sky130_fd_sc_hd__or3_1
X$13649 VPWR VGND VPWR \$1489 \$1462 VGND sky130_fd_sc_hd__inv_2
X$13650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13651 VGND \$1475 \$1034 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13652 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13653 VPWR \$1478 VPWR VGND \$1462 \$1477 \$1453 VGND sky130_fd_sc_hd__or3_1
X$13654 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13655 VGND \$1476 \$1248 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_8
X$13656 VGND \$1478 \$1490 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$13657 VGND \$1463 \$1342 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$13658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13660 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13661 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13664 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13665 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13666 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13667 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13668 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13670 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13671 VPWR \$1445 VGND VPWR \$1466 \$1342 VGND sky130_fd_sc_hd__or2_4
X$13672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13673 VPWR \$1454 VGND VPWR \$1219 \$1342 VGND sky130_fd_sc_hd__or2_4
X$13674 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13675 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13677 VPWR \$1425 VGND VPWR \$1058 \$1248 VGND sky130_fd_sc_hd__or2_4
X$13678 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13680 VPWR \$1342 VGND VPWR \$744 \$1434 VGND sky130_fd_sc_hd__or2_4
X$13681 VPWR \$1490 VGND VPWR \$1060 \$1401 VGND sky130_fd_sc_hd__or2_4
X$13682 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13684 VPWR \$1490 VGND VPWR \$1507 \$1425 VGND sky130_fd_sc_hd__or2_4
X$13685 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13686 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13687 VPWR \$1401 VGND VPWR \$433 \$1034 VGND sky130_fd_sc_hd__or2_4
X$13688 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13689 VPWR \$304 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13690 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13691 VPWR \$1508 \$304 VPWR \$1505 VGND \$1554 \$560 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$13692 VPWR \$1454 VGND VPWR \$325 \$1248 VGND sky130_fd_sc_hd__or2_4
X$13693 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13694 VPWR \$1490 VGND VPWR \$1421 \$1257 VGND sky130_fd_sc_hd__or2_4
X$13695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13696 VPWR \$1464 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13697 VGND \$1380 \$318 \$1464 \$1465 \$1266 \$601 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$13698 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13699 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13700 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13701 VGND \$1152 \$1455 \$605 \$1491 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13703 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13704 VPWR VGND \$1178 \$281 \$1455 \$1491 \$1166 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13705 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13706 VGND \$1152 \$1467 \$771 \$1479 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13707 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13708 VPWR VGND \$1178 \$200 \$1467 \$1479 \$1166 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13712 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13713 VPWR VPWR VGND \$1468 \$966 VGND sky130_fd_sc_hd__clkbuf_2
X$13714 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13715 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13716 VGND \$1152 \$1518 \$1203 \$1456 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13717 VGND \$1542 \$1202 \$1421 \$848 \$1155 \$1509 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$13718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13719 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13720 VGND \$1469 \$1480 \$1300 \$420 \$498 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$13721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13723 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13724 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13727 VGND \$358 \$1203 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$13728 VPWR VGND VPWR \$1480 \$1422 VGND sky130_fd_sc_hd__inv_2
X$13729 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13730 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13731 VPWR VGND \$1447 \$1644 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13733 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13734 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13735 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13737 VPWR \$1481 \$1413 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13738 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13740 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13741 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13742 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13744 VGND \$1152 \$1705 \$541 \$1492 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_4
X$13745 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13746 VGND \$1492 \$1705 \$1470 \$1222 \$2670 \$1011 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$13747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13749 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13750 VGND \$1152 \$1574 \$541 \$1510 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$13751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13752 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13753 VPWR VGND VPWR \$1470 \$1205 VGND sky130_fd_sc_hd__inv_2
X$13754 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13755 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13756 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13757 VPWR VGND VPWR \$1493 \$1520 VGND sky130_fd_sc_hd__inv_2
X$13758 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13759 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13760 VGND \$516 \$1576 \$541 \$1493 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13764 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13766 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13767 VPWR \$1511 VGND VPWR \$1494 \$1363 \$1482 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$13768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13769 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13770 VGND \$1494 \$1171 \$1450 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13772 VPWR VGND \$1311 \$1171 \$1450 \$1439 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13773 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13774 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13777 VGND \$516 \$1512 \$1274 \$1495 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13778 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13779 VGND \$1483 \$542 \$1430 \$1335 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13780 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13781 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13782 VPWR \$1495 VGND VPWR \$1483 \$1363 \$1512 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$13783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13784 VPWR \$1457 VGND VPWR \$1471 VGND sky130_fd_sc_hd__clkbuf_1
X$13785 VPWR VGND mgmt_gpio_oeb[3] VPWR \$1457 VGND sky130_fd_sc_hd__buf_2
X$13786 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13791 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13792 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13793 VPWR \$1028 \$853 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13794 VPWR VGND \$953 \$977 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13795 VPWR \$1039 VGND VPWR sram_ro_data[7] VGND sky130_fd_sc_hd__clkbuf_1
X$13796 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13799 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13800 VPWR VGND VPWR \$935 \$945 VGND sky130_fd_sc_hd__inv_2
X$13801 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13802 VPWR \$999 VGND \$945 VPWR \$906 VGND sky130_fd_sc_hd__nor2_1
X$13803 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13804 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13805 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13806 VPWR VGND \$564 \$790 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13807 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13808 VPWR \$639 VPWR VGND \$564 \$1014 \$1015 VGND sky130_fd_sc_hd__or3_1
X$13809 VPWR VGND VPWR \$428 \$639 VGND sky130_fd_sc_hd__inv_2
X$13810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13811 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13812 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13816 VPWR \$1041 VGND VPWR \$1029 VGND sky130_fd_sc_hd__clkbuf_1
X$13817 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13818 VPWR \$1029 VGND VPWR \$565 VGND sky130_fd_sc_hd__clkbuf_1
X$13819 VGND \$1016 \$1042 \$585 \$1014 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13820 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13821 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13822 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13823 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13824 VGND \$1001 \$986 \$381 \$1043 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$13825 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13826 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13828 VPWR \$1000 \$986 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13829 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13830 VPWR \$1001 VGND VPWR \$956 VGND sky130_fd_sc_hd__clkbuf_1
X$13831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13832 VGND \$987 \$1002 \$381 \$978 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$13833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13834 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13835 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13837 VPWR \$987 VGND VPWR \$957 VGND sky130_fd_sc_hd__clkbuf_1
X$13838 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13840 VGND \$308 \$1018 \$573 \$1045 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$13841 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13842 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13843 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13845 VPWR \$936 \$343 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13846 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13847 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13850 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13851 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13853 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13854 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13855 VGND \$856 \$979 \$922 \$1003 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13856 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13857 VPWR VGND \$701 \$293 \$979 \$1003 \$711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13858 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13859 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13860 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13861 VPWR VPWR VGND \$1032 \$711 VGND sky130_fd_sc_hd__clkbuf_2
X$13862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13863 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13864 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13865 VPWR VGND VPWR \$1004 \$959 VGND sky130_fd_sc_hd__inv_2
X$13866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13867 VPWR VGND \$792 \$200 \$980 \$960 \$793 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13868 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13869 VPWR VGND \$792 \$183 \$1005 \$989 \$793 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13870 VGND \$655 \$1005 \$961 \$989 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13871 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13872 VGND \$655 \$980 \$961 \$960 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13875 VGND \$463 \$961 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$13876 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13877 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13878 VPWR VGND \$892 \$281 \$981 \$1006 \$911 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13879 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13880 VPWR \$1007 \$939 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13883 VGND \$655 \$963 \$961 \$962 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13884 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13885 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13887 VPWR VPWR VGND \$1033 \$674 VGND sky130_fd_sc_hd__clkbuf_2
X$13888 VPWR VGND VPWR \$1019 \$963 VGND sky130_fd_sc_hd__inv_2
X$13889 VGND \$655 \$1061 \$605 \$1021 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$13890 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13891 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13892 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13893 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13894 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13897 VGND \$432 \$1034 \$1257 \$1022 \$1089 \$4275 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$13898 VGND \$463 \$605 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$13899 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13900 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13901 VGND \$900 \$1023 VPWR VPWR VGND sky130_fd_sc_hd__inv_8
X$13902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13903 VPWR \$964 VGND VPWR \$988 \$923 \$508 \$319 VGND
+ sky130_fd_sc_hd__o22a_1
X$13904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13905 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13906 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13908 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13909 VPWR \$1024 \$947 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$13910 VPWR VGND \$990 \$183 \$947 \$965 \$991 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13911 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13912 VPWR VGND \$990 \$294 \$1035 \$1062 \$991 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13914 VPWR VGND VPWR \$990 \$991 VGND sky130_fd_sc_hd__inv_2
X$13915 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13917 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13918 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13919 VPWR \$1025 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13920 VPWR \$992 VGND VPWR \$1025 VGND sky130_fd_sc_hd__clkbuf_1
X$13921 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13922 VGND \$1008 \$870 \$992 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13923 VPWR VGND \$713 \$200 \$949 \$967 \$714 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13925 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13926 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13927 VPWR \$3437 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13928 VGND \$1009 \$730 \$3437 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13929 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13930 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13932 VGND \$941 \$894 \$968 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13933 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13934 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13935 VPWR VGND \$713 \$184 \$982 \$994 \$714 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$13936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13937 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13938 VGND \$516 \$950 \$993 \$969 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13939 VGND \$516 \$982 \$993 \$994 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13940 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13941 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13943 VPWR \$1048 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13944 VGND \$951 \$950 \$1048 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13945 VGND \$872 \$982 \$983 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13946 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13947 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13948 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13949 VGND \$516 \$970 \$466 \$1010 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13950 VPWR \$1036 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13951 VPWR \$1036 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$13952 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13953 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13954 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13955 VGND \$1010 \$289 \$970 \$1026 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$13956 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13957 VGND \$516 \$1049 \$466 \$971 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13958 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13959 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13960 VGND \$942 \$952 \$1009 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$13961 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13963 VGND \$972 \$289 \$973 \$952 \$995 \$1027 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$13964 VPWR VGND VPWR \$1027 \$1008 VGND sky130_fd_sc_hd__inv_2
X$13965 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13966 VPWR VGND VPWR \$289 \$995 VGND sky130_fd_sc_hd__inv_4
X$13967 VGND \$516 \$974 \$466 \$996 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$13968 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13969 VGND \$996 \$289 \$973 \$974 \$1038 \$1037 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$13970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13971 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$13974 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13976 VPWR VGND \$895 \$1011 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$13977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13978 VGND \$1012 \$932 \$745 \$984 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$13979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13980 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13981 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13982 VGND \$1013 \$322 \$745 \$1011 \$934 \$975 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$13983 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13984 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$13985 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$13986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$13987 VPWR VGND VPWR \$943 \$997 VGND sky130_fd_sc_hd__inv_2
X$13988 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$13989 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$13990 VPWR \$984 VPWR VGND \$759 \$944 \$997 VGND sky130_fd_sc_hd__or3_1
X$13991 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13992 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$13993 VPWR VGND mgmt_gpio_out[1] VPWR \$1045 VGND sky130_fd_sc_hd__buf_2
X$13994 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13995 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13996 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13997 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$13998 VGND \$4093 \$4073 \$3531 \$3547 \$2221 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$13999 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14000 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14001 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14002 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14003 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14004 VPWR \$3994 VGND \$1963 \$2336 VPWR VGND sky130_fd_sc_hd__or2_1
X$14005 VPWR \$2815 \$3956 \$4074 \$3833 VGND \$3994 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$14006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14007 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14008 VPWR VGND VPWR \$4049 \$4075 VGND sky130_fd_sc_hd__inv_2
X$14009 VPWR VGND VPWR \$3472 \$4076 VGND sky130_fd_sc_hd__inv_2
X$14010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14011 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14012 VPWR \$4022 VGND \$4044 \$4061 VPWR VGND sky130_fd_sc_hd__or2_1
X$14013 VPWR \$3360 VGND \$4077 \$4061 VPWR VGND sky130_fd_sc_hd__or2_1
X$14014 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14015 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14016 VPWR \$4063 VGND \$4062 \$4078 VPWR VGND sky130_fd_sc_hd__or2_1
X$14017 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14018 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14019 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14023 VPWR \$3500 \$4095 \$2945 VPWR VGND \$4079 \$4080 VGND
+ sky130_fd_sc_hd__or4_1
X$14024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14025 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14027 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14028 VPWR \$3551 \$4012 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14029 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14030 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14031 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14032 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14033 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14034 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14035 VPWR VGND \$3894 \$4023 \$3998 \$4051 \$3908 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14036 VPWR VGND \$3894 \$281 \$4064 \$4096 \$3908 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14037 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14039 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14040 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14042 VGND \$4081 \$2539 \$2809 \$3218 \$2516 \$2295 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$14043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14044 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14045 VPWR \$4065 VGND VPWR \$3643 \$2254 \$4082 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$14046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14050 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14051 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14052 VPWR \$3535 VGND VPWR \$4053 \$1845 \$3963 \$1810 VGND
+ sky130_fd_sc_hd__o22a_1
X$14053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14054 VGND \$4083 \$4066 \$3162 \$2830 \$2651 \$3623 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14055 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14056 VPWR VGND VPWR \$3397 \$4083 \$4068 \$4067 \$4098 VGND
+ sky130_fd_sc_hd__and4_1
X$14057 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14058 VGND \$4067 \$4084 \$3936 \$2750 \$2541 \$3768 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14060 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14061 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14062 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14063 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14064 VPWR \$4099 VGND VPWR \$3923 \$2789 \$4085 \$1645 VGND
+ sky130_fd_sc_hd__o22a_1
X$14065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14066 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14067 VPWR \$4054 VGND VPWR \$2089 \$2559 \$4085 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$14068 VPWR VPWR VGND \$3769 \$4783 VGND sky130_fd_sc_hd__clkbuf_2
X$14069 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14070 VGND \$4016 \$4056 \$4085 \$2809 \$3218 \$4241 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14071 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14072 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14073 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14074 VPWR \$4100 VGND VPWR \$4086 \$2559 \$3402 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$14075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14076 VGND \$4101 \$4057 \$3825 \$2830 \$2651 \$1856 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14077 VGND \$3946 \$4059 \$3402 \$2809 \$3218 \$4087 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14079 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14080 VPWR \$1557 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14081 VPWR \$4069 VGND VPWR \$4088 \$2927 \$1557 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$14082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14083 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14087 VPWR \$4127 VGND \$2581 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$14088 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14089 VPWR \$3090 \$4089 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14090 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14091 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14092 VPWR \$3768 \$4090 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14094 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14095 VGND \$2989 \$4103 \$3590 \$4070 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14096 VPWR VGND VPWR \$3519 \$4091 VGND sky130_fd_sc_hd__inv_2
X$14097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14098 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14099 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14100 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14102 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14103 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14104 VPWR \$4071 VGND VPWR \$4092 VGND sky130_fd_sc_hd__clkbuf_1
X$14105 VPWR VGND mgmt_gpio_oeb[11] VPWR \$4071 VGND sky130_fd_sc_hd__buf_2
X$14106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14108 VGND \$4073 \$3277 \$4093 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$14109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14111 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14112 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14113 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14114 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14115 VPWR VGND VPWR \$3471 \$4113 VGND sky130_fd_sc_hd__inv_2
X$14116 VPWR VPWR \$4075 \$3880 VGND \$3742 VGND sky130_fd_sc_hd__nand2_2
X$14117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14118 VPWR \$3880 VPWR VGND \$4061 \$4062 VGND sky130_fd_sc_hd__or2_2
X$14119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14122 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14123 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14126 VPWR \$3011 \$4094 \$4010 VPWR VGND \$4129 \$4114 VGND
+ sky130_fd_sc_hd__or4_1
X$14127 VPWR \$4115 VGND \$4105 \$4130 \$2979 VPWR \$3492 VGND
+ sky130_fd_sc_hd__nor4_1
X$14128 VPWR VPWR VGND \$3126 \$4106 VGND sky130_fd_sc_hd__clkbuf_2
X$14129 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14130 VPWR \$4181 \$3838 \$4132 VPWR VGND \$4158 \$4080 VGND
+ sky130_fd_sc_hd__or4_1
X$14131 VPWR VGND VPWR \$4133 \$4131 VGND sky130_fd_sc_hd__inv_2
X$14132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14135 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14136 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14137 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14138 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14142 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14143 VGND \$856 \$4064 \$3921 \$4096 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14146 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14147 VPWR \$4081 VGND VPWR \$3814 \$2254 \$3898 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$14148 VGND \$3418 \$4116 \$3575 \$2809 \$3218 \$3537 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14149 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14150 VGND \$4065 \$2611 \$2809 \$3218 \$2477 \$2109 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$14151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14152 VPWR \$4097 VGND VPWR \$4117 \$2927 \$3364 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$14153 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14154 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14156 VPWR \$1235 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14157 VPWR \$4066 VGND VPWR \$4118 \$2927 \$1235 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$14158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14160 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14161 VGND \$4098 \$3938 \$2763 \$2369 \$2357 \$4119 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14162 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14163 VPWR \$4084 VGND VPWR \$4120 \$2559 \$1671 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$14164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14167 VGND \$3290 \$4099 \$4107 \$1625 \$1089 \$4134 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14170 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14171 VGND \$4015 \$4121 \$910 \$2525 \$2458 \$3748 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14173 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14174 VGND \$3900 \$4086 \$2031 \$1763 \$4122 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$14175 VGND \$4108 \$3985 \$4123 \$2369 \$2357 \$4293 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14176 VGND \$4125 \$4100 \$4124 \$2750 \$2541 \$3090 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14177 VPWR VGND VPWR \$4109 \$4101 \$4126 \$4125 \$4108 VGND
+ sky130_fd_sc_hd__and4_1
X$14178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14179 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14181 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14185 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14186 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14188 VPWR \$4135 VGND \$1645 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$14189 VPWR VGND \$3631 VPWR \$4127 VGND sky130_fd_sc_hd__clkbuf_4
X$14190 VPWR VGND \$3630 \$411 \$4089 \$4111 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14192 VPWR VGND \$3630 \$1171 \$4090 \$4102 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14193 VGND \$2989 \$4090 \$3590 \$4102 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$14194 VPWR VGND \$3716 \$386 \$4103 \$4070 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14195 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14197 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14198 VPWR VGND \$3716 \$542 \$4128 \$4136 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14200 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14201 VPWR VGND VPWR \$3872 \$3851 VGND sky130_fd_sc_hd__inv_2
X$14202 VGND \$2989 \$4190 \$3590 \$4112 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14203 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14204 VPWR \$4092 VGND VPWR \$2671 VGND sky130_fd_sc_hd__clkbuf_1
X$14205 VPWR \$4110 \$3010 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14206 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14208 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14210 VPWR VGND wb_dat_o[20] VPWR \$4949 VGND sky130_fd_sc_hd__buf_2
X$14211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14212 VPWR \$4976 VGND VPWR \$4950 \$4508 \$1769 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$14213 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14216 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14217 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14218 VPWR \$4864 \$4908 \$4733 VPWR VGND \$4891 \$4880 VGND
+ sky130_fd_sc_hd__or4_1
X$14219 VPWR \$4833 \$4929 \$4733 VPWR VGND \$4891 \$4880 VGND
+ sky130_fd_sc_hd__or4_1
X$14220 VPWR VGND \$3833 VPWR \$4929 VGND sky130_fd_sc_hd__clkbuf_4
X$14221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14223 VPWR \$4909 VPWR VGND \$4930 \$4942 \$3742 VGND sky130_fd_sc_hd__or3b_1
X$14224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14225 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14226 VPWR \$4941 \$4917 VGND \$4930 VPWR \$4212 \$4698 VGND
+ sky130_fd_sc_hd__or4_2
X$14227 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14228 VGND \$4951 \$2815 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$14229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14230 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14231 VGND \$4733 \$3155 \$4833 \$4853 \$4891 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$14232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14233 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14234 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14235 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14236 VGND \$4568 \$4931 \$4930 \$4735 \$4664 \$5040 VPWR VPWR VGND
+ sky130_fd_sc_hd__a41o_1
X$14237 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14238 VPWR \$4735 VGND \$4918 \$4855 VPWR VGND sky130_fd_sc_hd__or2_1
X$14239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14242 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14243 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14244 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14245 VPWR VGND \$4912 VPWR \$2640 \$4952 \$4962 VGND sky130_fd_sc_hd__a21oi_1
X$14246 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14249 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14250 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14251 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14252 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14253 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14254 VPWR \$4739 VGND \$2815 VPWR \$4953 VGND sky130_fd_sc_hd__nor2_1
X$14255 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14256 VGND \$4952 \$4963 \$4665 \$4758 VPWR VPWR \$4739 VGND
+ sky130_fd_sc_hd__or4b_1
X$14257 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14258 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14259 VPWR \$4605 VGND \$4964 \$4954 VPWR VGND sky130_fd_sc_hd__or2_1
X$14260 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14261 VPWR \$4580 VPWR VGND \$4954 \$4913 \$4932 VGND sky130_fd_sc_hd__or3_1
X$14262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14264 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14265 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14267 VPWR \$1725 \$1712 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$14268 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14269 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14270 VPWR \$1725 VPWR \$4933 VGND \$4934 \$4897 \$4921 VGND
+ sky130_fd_sc_hd__o211a_2
X$14271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14272 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14273 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14274 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14275 VGND \$2777 \$4923 \$4811 \$4922 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14276 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14277 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14280 VPWR VGND VPWR \$4760 \$4717 VGND sky130_fd_sc_hd__inv_2
X$14281 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14282 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14283 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14284 VGND \$4761 \$4935 \$4811 \$4943 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14285 VPWR VGND \$4760 \$4023 \$4935 \$4943 \$4717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14286 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14287 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14288 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14289 VPWR VGND \$4955 \$2516 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$14290 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14291 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14292 VPWR VGND \$4935 \$2477 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$14293 VPWR VGND \$4781 \$3732 \$4944 \$4965 \$4782 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14294 VPWR VGND VPWR \$4781 \$4782 VGND sky130_fd_sc_hd__inv_2
X$14295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14296 VPWR VGND \$4781 \$4023 \$4967 \$4966 \$4782 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14297 VPWR VGND VPWR \$2783 \$4944 VGND sky130_fd_sc_hd__inv_2
X$14298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14299 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14300 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14301 VPWR VGND VPWR \$2611 \$4967 VGND sky130_fd_sc_hd__inv_2
X$14302 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14303 VGND \$4761 \$4936 \$4813 \$4956 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$14304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14305 VPWR VGND \$4654 \$542 \$4936 \$4956 \$4667 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14306 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14307 VGND \$3037 \$4936 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$14308 VGND \$4761 \$4937 \$4813 \$4968 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14309 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14310 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14311 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14312 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14313 VPWR VGND VPWR \$3405 \$4937 VGND sky130_fd_sc_hd__inv_2
X$14314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14316 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14317 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14319 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14320 VPWR VGND \$5005 \$1179 \$4958 \$4969 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14321 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14322 VPWR \$4945 VGND \$2375 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$14323 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14324 VPWR VGND \$4957 VPWR \$4945 VGND sky130_fd_sc_hd__clkbuf_4
X$14325 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14326 VPWR \$3965 \$4958 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14328 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14329 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14331 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14332 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14333 VPWR \$3645 \$4959 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14335 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14336 VPWR VGND \$4905 \$1179 \$4959 \$4970 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14337 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14338 VGND \$4764 \$4901 \$4850 \$4914 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14341 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14342 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14343 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14344 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14345 VPWR VGND VPWR \$2531 \$4982 VGND sky130_fd_sc_hd__inv_2
X$14346 VGND \$4764 \$4938 \$4765 \$4971 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14347 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14348 VPWR \$3944 \$4938 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14351 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14352 VPWR \$3095 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14353 VGND \$3438 \$4481 \$3095 \$4926 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$14354 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14355 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14356 VPWR VGND \$4899 \$542 \$4960 \$4972 \$4900 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14357 VPWR VGND VPWR \$4481 \$4960 VGND sky130_fd_sc_hd__inv_2
X$14358 VPWR VGND VPWR \$4899 \$4900 VGND sky130_fd_sc_hd__inv_2
X$14359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14360 VPWR \$4973 VGND \$2614 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$14361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14363 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14364 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14367 VGND \$4764 \$4925 \$5006 \$4924 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14371 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14374 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14375 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14377 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14378 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14379 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14380 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14383 VPWR \$4961 VGND VPWR \$4946 VGND sky130_fd_sc_hd__clkbuf_1
X$14384 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14385 VGND \$4946 \$4939 \$386 \$4686 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$14386 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14387 VGND \$2989 \$4939 \$4828 \$4961 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$14388 VPWR VGND \$4939 \$3107 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$14389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14390 VGND \$4948 \$5034 \$4974 \$4939 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$14391 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14392 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14395 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14396 VGND \$2989 \$4940 \$4828 \$4947 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14397 VPWR VGND \$4650 \$386 \$4940 \$4947 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14399 VGND \$4878 \$386 \$4940 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$14400 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14401 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14402 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14403 VGND \$4948 mgmt_gpio_out[14] \$3036 VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_2
X$14404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14406 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14407 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14408 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14409 VPWR debug_out VPWR VGND \$839 VGND sky130_fd_sc_hd__buf_4
X$14410 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14415 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14418 VPWR \$2698 VGND \$2659 \$2552 VPWR VGND sky130_fd_sc_hd__or2_1
X$14419 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14420 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14421 VGND \$2713 \$2740 \$2741 \$2659 \$2659 \$2700 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14422 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14423 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14425 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14426 VPWR \$2758 VGND \$2514 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$14427 VPWR VGND VPWR \$2795 \$2758 VGND sky130_fd_sc_hd__inv_2
X$14428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14429 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14430 VPWR \$2714 VGND \$2453 VPWR \$2742 VGND sky130_fd_sc_hd__nor2_1
X$14431 VPWR \$2743 VGND \$2714 VPWR \$2679 VGND sky130_fd_sc_hd__nor2_1
X$14432 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14434 VPWR \$2744 VGND \$2453 \$2815 VPWR VGND sky130_fd_sc_hd__or2_1
X$14435 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14436 VPWR \$2743 \$2701 VPWR \$2744 VGND VGND sky130_fd_sc_hd__and2_1
X$14437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14439 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14440 VPWR \$2796 VGND \$2392 \$2745 VPWR VGND sky130_fd_sc_hd__or2_1
X$14441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14442 VPWR \$2745 VGND \$2488 VPWR \$2815 VGND sky130_fd_sc_hd__nor2_1
X$14443 VPWR \$2731 VGND \$2745 VPWR \$2717 VGND sky130_fd_sc_hd__nor2_1
X$14444 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14445 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14446 VPWR VPWR \$2741 VGND \$2488 \$2759 \$2746 VGND sky130_fd_sc_hd__o21ai_1
X$14447 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14448 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14449 VPWR \$2488 VPWR \$2746 VGND \$2731 \$2700 VGND sky130_fd_sc_hd__o21a_1
X$14450 VPWR \$2797 VGND \$2553 \$2774 VPWR VGND sky130_fd_sc_hd__or2_1
X$14451 VPWR VGND \$2741 \$2640 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$14452 VGND \$856 \$2702 \$1750 \$2760 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14453 VPWR \$2798 VGND \$2774 VPWR \$2759 VGND sky130_fd_sc_hd__nor2_1
X$14454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14455 VPWR VGND \$2775 \$293 \$2702 \$2760 \$2776 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14456 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14458 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14459 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14460 VPWR VGND \$2775 \$294 \$2732 \$2761 \$2776 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14461 VGND \$856 \$2732 \$2556 \$2761 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14463 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14464 VGND \$856 \$2733 \$1861 \$2762 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$14465 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14466 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14467 VGND \$856 \$2777 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$14468 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14469 VGND \$2762 \$1183 \$183 \$2778 \$2779 \$2733 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14470 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14472 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14473 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14475 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14476 VGND \$856 \$2764 \$2556 \$2799 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14477 VGND \$856 \$2704 \$2556 \$2718 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14478 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14479 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14481 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14482 VPWR \$1490 VGND VPWR \$2734 \$1444 VGND sky130_fd_sc_hd__or2_4
X$14483 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14484 VPWR \$2800 VGND VPWR \$2719 \$1954 \$2780 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$14485 VPWR \$2123 \$2764 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14486 VGND \$2782 \$2575 \$2749 \$1065 \$880 \$2781 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14487 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14488 VPWR \$2735 VGND VPWR \$2747 \$2456 \$2748 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$14489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14490 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14492 VPWR VGND VPWR \$2802 \$2765 \$2801 \$2782 \$2328 VGND
+ sky130_fd_sc_hd__and4_1
X$14493 VGND \$2765 \$2686 \$769 \$2073 \$2096 \$2748 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14494 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14495 VPWR \$2766 VGND VPWR \$769 \$2559 \$2783 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$14496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14498 VGND \$2722 \$2720 \$495 \$2369 \$2357 \$2749 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14500 VGND \$2723 \$2766 \$2780 \$2750 \$2541 \$796 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14501 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14503 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14504 VPWR \$2767 VGND VPWR \$1072 \$686 \$2763 \$1466 VGND
+ sky130_fd_sc_hd__o22a_1
X$14505 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14506 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14507 VGND \$1765 \$2767 \$2383 \$2372 \$2497 \$2784 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14511 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14512 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14513 VPWR \$1570 VGND VPWR \$2785 \$1264 VGND sky130_fd_sc_hd__or2_4
X$14514 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14515 VPWR \$1570 VGND VPWR \$2751 \$1283 VGND sky130_fd_sc_hd__or2_4
X$14516 VGND \$2786 \$2612 \$2804 \$2162 \$2384 \$2123 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14517 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14518 VPWR VGND VPWR \$1624 \$2786 \$2803 \$449 \$2787 VGND
+ sky130_fd_sc_hd__and4_1
X$14519 VPWR \$2768 VGND VPWR \$2749 \$2366 \$1240 \$1558 VGND
+ sky130_fd_sc_hd__o22a_1
X$14520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14522 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14523 VGND \$2769 \$2788 \$2747 \$1340 \$1625 \$2753 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14524 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14525 VGND \$2726 \$754 \$2752 \$2789 \$2372 \$2719 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14526 VGND \$2805 \$1696 \$2790 \$2789 \$1507 \$756 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14529 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14530 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14532 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14534 VGND \$2807 \$2768 \$2503 \$2785 \$2751 \$2691 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14535 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14536 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14537 VPWR \$2728 VGND VPWR \$2561 \$2665 \$2753 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$14538 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14539 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14540 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14541 VPWR VPWR VGND \$2808 \$1468 VGND sky130_fd_sc_hd__clkbuf_2
X$14542 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14545 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14546 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14548 VPWR \$2770 VGND VPWR \$2923 \$2559 \$1892 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$14549 VGND \$2792 \$2770 \$1821 \$2750 \$2541 \$2791 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14550 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14551 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14552 VPWR VGND VPWR \$2754 \$2811 \$2810 \$2792 \$2793 VGND
+ sky130_fd_sc_hd__and4_1
X$14553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14554 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14555 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14557 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14559 VGND \$2771 \$2794 \$1521 \$2665 \$2688 \$2111 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14560 VGND \$2754 \$2771 \$2755 \$2692 VPWR \$1048 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$14561 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14562 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14563 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14565 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14566 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14567 VGND \$2812 \$2772 \$2033 \$2047 \$2048 \$2791 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14568 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14569 VPWR \$2772 VGND VPWR \$2403 \$1956 \$1225 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$14570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14572 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14573 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14576 VGND \$1152 \$2709 \$2450 \$2736 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14578 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14580 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14581 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14582 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14583 VPWR VGND \$2653 \$1927 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$14584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14586 VPWR VGND \$2694 \$542 \$2729 \$2737 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14587 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14588 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14590 VGND \$1152 \$2729 \$2450 \$2737 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14591 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14592 VPWR \$2813 \$2773 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14593 VPWR VGND \$2730 \$411 \$2773 \$2738 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14594 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14595 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14596 VGND \$1152 \$2773 \$2232 \$2738 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14597 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14598 VPWR \$2730 \$2711 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14600 VPWR VGND \$2730 \$542 \$2696 \$2673 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14602 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14603 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14604 VPWR \$2739 VGND VPWR mgmt_gpio_in[7] VGND sky130_fd_sc_hd__clkbuf_1
X$14605 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14606 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14607 VPWR VGND VPWR \$2739 \$2756 VGND sky130_fd_sc_hd__inv_4
X$14608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14609 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14610 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14611 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14612 VPWR VGND \$5877 VPWR wb_stb_i VGND sky130_fd_sc_hd__clkbuf_4
X$14613 VPWR VGND wb_ack_o VPWR \$3831 VGND sky130_fd_sc_hd__buf_2
X$14614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14615 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14617 VPWR VPWR \$3470 VGND \$2320 \$3852 \$3853 VGND sky130_fd_sc_hd__o21ai_1
X$14618 VPWR VGND \$3832 \$3852 \$3409 VPWR \$3097 \$3805 VGND
+ sky130_fd_sc_hd__or4b_2
X$14619 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14620 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14621 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14622 VPWR \$3853 VPWR VGND \$2234 \$3470 VGND sky130_fd_sc_hd__or2_2
X$14623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14624 VPWR \$3661 VGND \$2119 VPWR \$3833 VGND sky130_fd_sc_hd__nor2_1
X$14625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14626 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14628 VPWR VGND VPWR \$3855 \$3758 VGND sky130_fd_sc_hd__inv_2
X$14629 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14630 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14631 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14632 VPWR \$3855 \$3257 VGND \$3681 VPWR \$3806 \$3834 VGND
+ sky130_fd_sc_hd__or4_2
X$14633 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14634 VPWR \$3834 VGND \$3878 \$3689 VPWR VGND sky130_fd_sc_hd__or2_1
X$14635 VPWR \$3775 VPWR VGND \$3855 \$3856 \$3834 VGND sky130_fd_sc_hd__or3_1
X$14636 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14637 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14638 VPWR VGND VPWR \$3879 \$3502 VGND sky130_fd_sc_hd__inv_2
X$14639 VGND \$3742 \$3491 \$3835 \$3836 \$3124 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22ai_2
X$14640 VGND \$3835 \$3879 \$3862 \$3880 \$3742 \$3836 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_4
X$14641 VPWR \$3835 VGND \$3501 VPWR \$3857 VGND sky130_fd_sc_hd__nor2_1
X$14642 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14643 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14644 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14645 VGND \$3473 \$3452 \$3472 \$3858 \$3779 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$14646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14649 VPWR \$3777 VPWR VGND \$3788 \$3789 \$3859 VGND sky130_fd_sc_hd__or3b_1
X$14650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14651 VPWR \$2741 \$3788 \$2949 \$2996 VGND \$3709 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$14652 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14653 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14654 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14655 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14657 VPWR \$3789 \$3861 \$3343 VPWR VGND \$3860 \$3474 VGND
+ sky130_fd_sc_hd__or4_1
X$14658 VPWR \$3881 VGND \$3710 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$14659 VPWR VGND VPWR \$3789 \$3881 VGND sky130_fd_sc_hd__inv_2
X$14660 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14661 VPWR \$4010 \$3793 \$3861 VPWR VGND \$2979 \$2945 VGND
+ sky130_fd_sc_hd__or4_1
X$14662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14663 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14665 VGND \$3792 \$3862 \$2990 \$3500 \$3810 \$3837 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$14666 VPWR \$3874 VGND \$3759 VPWR \$3778 VGND sky130_fd_sc_hd__nor2_1
X$14667 VPWR \$3863 VGND \$3862 VPWR \$3793 VGND sky130_fd_sc_hd__nor2_1
X$14668 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14669 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14670 VPWR VGND VPWR \$3790 \$3882 VGND sky130_fd_sc_hd__inv_2
X$14671 VPWR \$3597 \$3561 VPWR \$3863 \$3838 \$3882 VGND \$3874 VGND
+ sky130_fd_sc_hd__o221ai_1
X$14672 VPWR VGND VPWR \$3837 \$3838 VGND sky130_fd_sc_hd__inv_2
X$14673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14674 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14675 VGND \$2777 \$3812 \$3413 \$3811 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$14676 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14678 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14679 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14680 VGND \$2777 \$3839 \$3413 \$3875 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14681 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14682 VPWR VGND VPWR \$3864 \$3812 VGND sky130_fd_sc_hd__inv_2
X$14683 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14684 VPWR VGND \$3670 \$293 \$3839 \$3875 \$3653 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14687 VPWR VGND VPWR \$2296 \$3839 VGND sky130_fd_sc_hd__inv_2
X$14688 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14690 VGND \$3732 \$294 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$14691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14693 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14694 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14695 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14697 VPWR \$2595 VGND VPWR \$3883 \$3562 \$2819 \$3621 VGND
+ sky130_fd_sc_hd__o22a_1
X$14698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14699 VPWR VGND VPWR \$2748 \$3884 VGND sky130_fd_sc_hd__inv_2
X$14700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14701 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14704 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14706 VPWR \$3865 VGND VPWR \$2539 \$3556 \$2281 \$3106 VGND
+ sky130_fd_sc_hd__o22a_1
X$14707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14710 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14711 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14713 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14714 VPWR \$3841 VGND VPWR \$1019 \$1060 \$3712 \$3703 VGND
+ sky130_fd_sc_hd__o22a_1
X$14715 VGND \$3797 \$3841 \$2515 \$3271 \$3019 \$3842 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14716 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14720 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14721 VGND \$3816 \$3865 \$3814 \$3562 \$3765 \$3796 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14722 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14723 VPWR \$1293 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14724 VPWR VGND VPWR \$3885 \$1293 VGND sky130_fd_sc_hd__inv_2
X$14725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14726 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14728 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14729 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14730 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14731 VPWR \$1466 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14732 VGND \$2582 \$3843 \$3935 \$1810 \$1466 \$3236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14733 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14734 VPWR \$3843 VGND VPWR \$3864 \$3042 \$3723 \$2447 VGND
+ sky130_fd_sc_hd__o22a_1
X$14735 VGND \$3819 \$3374 \$3886 \$2918 \$3181 \$3898 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14738 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14740 VGND \$3867 \$3844 \$2516 \$2734 \$2031 \$3866 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14742 VPWR VGND VPWR \$3781 \$3823 \$3845 \$3867 \$3868 VGND
+ sky130_fd_sc_hd__and4_1
X$14743 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14745 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14747 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14748 VPWR \$3869 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14749 VPWR \$3672 \$3870 VPWR \$3910 VGND \$3562 \$3869 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$14750 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14751 VPWR \$3870 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14752 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14753 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14754 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14755 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14757 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14758 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14759 VGND \$3871 \$3847 \$3846 \$3824 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$14760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14761 VPWR \$3846 VGND VPWR \$3541 \$3765 \$3090 \$2581 VGND
+ sky130_fd_sc_hd__o22a_1
X$14762 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14764 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14766 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14768 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14769 VGND \$3848 \$3826 \$3771 \$2750 \$2541 \$3628 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14770 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14771 VGND \$3850 \$3887 \$3828 \$2830 \$2651 \$3338 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14772 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14773 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14774 VPWR VGND VPWR \$3406 \$3850 \$3849 \$3848 \$3827 VGND
+ sky130_fd_sc_hd__and4_1
X$14775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14777 VGND \$3735 \$3772 \$2430 \$2809 \$3218 \$4279 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14778 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14780 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14781 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14783 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14784 VGND \$2989 \$3802 \$4164 \$3829 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14786 VPWR VGND VPWR \$3628 \$3802 VGND sky130_fd_sc_hd__inv_2
X$14787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14789 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14793 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14794 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14795 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14796 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14797 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14798 VGND \$2989 \$3888 \$3590 \$3876 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$14799 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14801 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14802 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14803 VPWR VGND \$3872 \$354 \$3803 \$3785 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14804 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14806 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14807 VPWR VGND \$3872 \$1179 \$3756 \$3877 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14808 VGND \$2989 \$3756 \$3590 \$3877 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$14809 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14810 VGND \$3889 \$780 \$3890 \$482 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$14811 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14812 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14813 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14814 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14815 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14816 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14818 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14819 VPWR VGND wb_dat_o[6] VPWR \$4264 VGND sky130_fd_sc_hd__buf_2
X$14820 VPWR \$4324 VGND VPWR \$4264 \$3531 \$1769 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$14821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14825 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14826 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14828 VPWR \$4034 VPWR VGND \$3498 \$3430 \$4299 VGND sky130_fd_sc_hd__or3_2
X$14829 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14830 VPWR VPWR \$3616 VGND \$4265 \$2214 \$4325 \$3648 VGND
+ sky130_fd_sc_hd__a211o_1
X$14831 VPWR VGND VPWR \$4325 \$4193 VGND sky130_fd_sc_hd__inv_2
X$14832 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14833 VPWR VPWR VGND \$4266 \$3277 VGND sky130_fd_sc_hd__clkbuf_2
X$14834 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14835 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14836 VPWR VGND \$2996 VPWR \$1998 \$4300 \$3470 VGND sky130_fd_sc_hd__a21oi_1
X$14837 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14838 VGND \$3759 \$4305 \$3856 \$3906 \$4410 \$4300 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2111o_2
X$14839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14840 VPWR \$4306 VPWR \$3995 VGND \$4138 \$4214 VGND sky130_fd_sc_hd__o21a_1
X$14841 VPWR VPWR \$4307 VGND \$4337 \$4138 \$4308 VGND sky130_fd_sc_hd__o21ai_1
X$14842 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14844 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14845 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14846 VPWR VGND VPWR \$4307 \$4215 VGND sky130_fd_sc_hd__inv_2
X$14847 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14850 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14851 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14852 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14853 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14855 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14856 VGND \$4253 \$2444 \$3255 \$4268 \$4267 VPWR VPWR VGND
+ sky130_fd_sc_hd__nor4_2
X$14857 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14858 VGND \$4301 \$3806 \$3260 \$4309 \$4326 VPWR VPWR VGND
+ sky130_fd_sc_hd__nor4_2
X$14859 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14860 VPWR \$4079 VPWR VGND \$4267 \$4286 \$4115 VGND sky130_fd_sc_hd__or3_1
X$14861 VPWR \$4115 VGND \$4310 VPWR \$3892 VGND sky130_fd_sc_hd__nor2_1
X$14862 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14863 VPWR \$4154 VGND \$4310 VPWR \$2815 VGND sky130_fd_sc_hd__nor2_1
X$14864 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14865 VGND \$4311 \$4156 \$3666 \$4253 \$4301 \$4312 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_4
X$14866 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14867 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14868 VPWR \$4094 \$4287 \$4131 VPWR VGND \$4154 \$4269 VGND
+ sky130_fd_sc_hd__or4_1
X$14869 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14870 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14872 VPWR VGND \$4234 \$3711 \$4254 \$4233 \$4224 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14873 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14874 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14875 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14876 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14877 VPWR VGND \$4234 \$293 \$4327 \$4328 \$4224 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14878 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14879 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14880 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14881 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14882 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14883 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14884 VPWR \$3712 \$4327 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$14885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14886 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14887 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14888 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14889 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14890 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14891 VGND \$2777 \$4271 \$3921 \$4288 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14892 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14893 VPWR VGND \$4270 \$3732 \$4271 \$4288 \$4272 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14894 VPWR \$4289 VGND \$2734 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$14895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14896 VPWR \$4290 VGND \$3271 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$14897 VPWR VPWR VGND \$4290 \$4272 VGND sky130_fd_sc_hd__clkbuf_2
X$14898 VPWR VGND VPWR \$2840 \$4271 VGND sky130_fd_sc_hd__inv_2
X$14899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14901 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14902 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14908 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14911 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14912 VPWR \$4329 VGND \$3271 \$2610 VPWR VGND sky130_fd_sc_hd__or2_1
X$14913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14915 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14916 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14919 VGND \$4313 \$4144 \$4314 \$4329 \$3019 \$4118 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$14920 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14921 VPWR \$4273 VGND VPWR \$1838 \$2456 \$4274 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$14922 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14923 VGND \$4068 \$4273 \$4275 \$2525 \$2458 \$3979 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14924 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14925 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14928 VGND \$4276 \$1118 \$4302 \$3818 VPWR VPWR VGND sky130_fd_sc_hd__and3_4
X$14929 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14930 VGND \$4330 \$3696 \$4120 \$2073 \$2096 \$4274 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14931 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$14933 VPWR \$4240 VGND VPWR \$3350 \$2456 \$4027 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$14934 VPWR \$4161 VGND VPWR \$4315 \$2447 \$3581 \$3765 VGND
+ sky130_fd_sc_hd__o22a_1
X$14935 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14936 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14938 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14939 VPWR \$4257 VGND VPWR \$910 \$2135 \$3399 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$14940 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14941 VGND \$4331 \$4257 \$3886 \$1065 \$880 \$2397 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14942 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14943 VGND \$4291 \$3376 \$3866 \$2073 \$2096 \$4145 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14944 VPWR \$4242 VGND VPWR \$4134 \$2135 \$2163 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$14945 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14946 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14947 VPWR \$929 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14948 VGND \$3770 \$4277 \$4292 VPWR \$929 VPWR VGND sky130_fd_sc_hd__nand3_4
X$14949 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14950 VPWR VGND VPWR \$4277 \$4291 \$4316 \$4331 \$4317 VGND
+ sky130_fd_sc_hd__and4_1
X$14951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14953 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14954 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14955 VPWR \$4318 VGND VPWR \$4278 \$2135 \$4319 \$2107 VGND
+ sky130_fd_sc_hd__o22a_1
X$14956 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14957 VPWR \$4122 VGND VPWR \$4258 \$1819 \$4124 \$1845 VGND
+ sky130_fd_sc_hd__o22a_1
X$14958 VGND \$4332 \$4318 \$4293 \$1065 \$880 \$3584 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14959 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14960 VGND \$4126 \$4259 \$4278 \$2525 \$2458 \$4087 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$14962 VGND \$4333 \$3273 \$4086 \$2073 \$2096 \$4243 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14963 VPWR \$3799 VGND VPWR \$4243 \$2986 \$4293 \$2918 VGND
+ sky130_fd_sc_hd__o22a_1
X$14964 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14965 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14966 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14967 VGND \$3947 \$4343 \$4417 VPWR \$862 VPWR VGND sky130_fd_sc_hd__nand3_4
X$14968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$14969 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14970 VPWR \$862 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$14971 VGND \$3849 \$4260 \$4294 \$2525 \$2458 \$4279 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14973 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14974 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14975 VGND \$4334 \$3380 \$3783 \$2073 \$2096 \$4244 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14976 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14978 VGND \$4296 \$4295 \$3112 \$1879 \$2031 \$4031 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14979 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14980 VPWR \$4335 VGND \$2031 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$14981 VGND \$4281 \$4320 \$3678 \$1561 \$3765 \$3929 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$14982 VPWR \$4280 \$4296 \$4281 VGND VPWR \$3224 VGND sky130_fd_sc_hd__and3_2
X$14983 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14984 VGND \$2989 \$4245 \$4164 \$4297 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14985 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14987 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14988 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14989 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14990 VGND \$2989 \$4189 \$4164 \$4346 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$14991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$14992 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$14993 VPWR \$4298 VGND \$3765 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$14994 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$14995 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$14996 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$14997 VPWR VGND VPWR \$4187 \$4282 VGND sky130_fd_sc_hd__inv_2
X$14998 VPWR VGND \$4303 \$184 \$4282 \$4336 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$14999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15000 VPWR \$3979 \$4283 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15001 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15002 VGND \$2989 \$4283 \$4165 \$4284 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15003 VPWR VGND \$4303 \$1171 \$4283 \$4284 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15005 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15006 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15007 VGND \$2989 \$4246 \$4165 \$4322 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15008 VGND \$3952 \$3633 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$15009 VPWR VGND \$3851 VPWR \$4298 VGND sky130_fd_sc_hd__clkbuf_4
X$15010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15011 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15013 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15014 VPWR VGND \$3872 \$184 \$4247 \$4262 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15015 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15016 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15017 VPWR VGND \$3872 \$542 \$4285 \$4348 \$3851 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15018 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15019 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15020 VGND \$2866 \$4285 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$15021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15023 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15024 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15025 VPWR \$4248 VGND VPWR mgmt_gpio_in[12] VGND sky130_fd_sc_hd__clkbuf_1
X$15026 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15028 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15029 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15030 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15031 VPWR \$1263 VGND VPWR sram_ro_data[11] VGND sky130_fd_sc_hd__clkbuf_1
X$15032 VPWR VGND VPWR \$1267 \$1263 VGND sky130_fd_sc_hd__inv_2
X$15033 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15034 VPWR \$1276 VGND VPWR sram_ro_data[12] VGND sky130_fd_sc_hd__clkbuf_1
X$15035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15036 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15037 VPWR \$1277 VGND VPWR \$1269 VGND sky130_fd_sc_hd__clkbuf_1
X$15038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15039 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15040 VPWR \$1278 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$15041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15043 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15045 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15046 VPWR VGND VPWR \$1042 \$1292 VGND sky130_fd_sc_hd__inv_2
X$15047 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15049 VPWR VGND VPWR \$1254 \$1187 VGND sky130_fd_sc_hd__inv_2
X$15050 VPWR \$1279 VGND \$1188 \$1042 VPWR VGND sky130_fd_sc_hd__or2_1
X$15051 VPWR VGND VPWR \$1188 \$1014 VGND sky130_fd_sc_hd__inv_2
X$15052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15053 VPWR \$1255 VPWR VGND \$564 \$1188 \$1015 VGND sky130_fd_sc_hd__or3_1
X$15054 VGND \$1255 \$1078 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$15055 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15056 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15057 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15058 VPWR \$1280 VGND VPWR \$1270 VGND sky130_fd_sc_hd__clkbuf_1
X$15059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15060 VGND \$1243 \$1215 \$387 \$1227 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$15061 VPWR \$1281 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$15062 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15063 VPWR \$1243 VGND VPWR \$1281 VGND sky130_fd_sc_hd__clkbuf_1
X$15064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15065 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15066 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15067 VPWR \$1245 VGND VPWR \$1228 VGND sky130_fd_sc_hd__clkbuf_1
X$15068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15069 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15071 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15072 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15073 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15076 VGND \$1230 \$780 \$986 \$1015 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$15077 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15079 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15081 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15082 VGND \$856 \$1231 \$891 \$1209 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15083 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15084 VGND \$655 \$856 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$15085 VPWR VGND VPWR \$1282 \$1231 VGND sky130_fd_sc_hd__inv_2
X$15086 VPWR VGND \$1146 \$1265 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$15087 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15088 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15089 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15090 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15092 VPWR VPWR VGND \$1246 \$1088 VGND sky130_fd_sc_hd__clkbuf_2
X$15093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15095 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15096 VPWR \$1256 \$1216 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15098 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15099 VPWR \$1246 VGND \$1271 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$15100 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15102 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15103 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15104 VGND \$1175 \$1233 \$183 \$1217 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$15105 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15107 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15108 VPWR VGND VPWR \$1232 \$1233 VGND sky130_fd_sc_hd__inv_2
X$15109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15110 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15111 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15113 VPWR \$1257 VGND VPWR \$1114 \$1248 VGND sky130_fd_sc_hd__or2_4
X$15114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15115 VPWR \$1218 VGND \$1258 \$1248 VPWR VGND sky130_fd_sc_hd__or2_1
X$15116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15118 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15120 VPWR VGND VPWR \$1259 \$1195 VGND sky130_fd_sc_hd__inv_2
X$15121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15122 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15123 VPWR \$566 VPWR VGND \$1264 \$1248 VGND sky130_fd_sc_hd__or2_2
X$15124 VPWR \$353 VPWR VGND \$1283 \$1034 VGND sky130_fd_sc_hd__or2_2
X$15125 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15131 VGND \$655 \$1293 \$605 \$1285 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$15132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15133 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15134 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15135 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15137 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15138 VPWR VGND VPWR \$1242 \$1177 VGND sky130_fd_sc_hd__inv_2
X$15139 VGND \$655 \$1250 \$605 \$1249 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15141 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15142 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15143 VGND \$1251 \$499 \$1221 \$1198 \$1266 \$684 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15146 VPWR VGND VPWR \$1178 \$1166 VGND sky130_fd_sc_hd__inv_2
X$15147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15150 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15152 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15153 VGND \$1152 \$1252 \$771 \$1272 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15154 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15155 VPWR VGND \$990 \$1179 \$1252 \$1272 \$991 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15157 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15159 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15160 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15161 VGND \$1152 \$1287 \$1203 \$1286 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15162 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15163 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15164 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15165 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15166 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15170 VPWR \$1253 VGND \$1198 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$15171 VPWR VGND \$1182 VPWR \$1253 VGND sky130_fd_sc_hd__clkbuf_4
X$15172 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15173 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15174 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15175 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15176 VPWR VGND VPWR \$1170 \$1182 VGND sky130_fd_sc_hd__inv_2
X$15177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15180 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15181 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15182 VGND \$358 \$993 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$15183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15184 VPWR VGND VPWR \$1260 \$1137 VGND sky130_fd_sc_hd__inv_2
X$15185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15188 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15190 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15191 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15192 VPWR VPWR VGND \$1066 \$541 VGND sky130_fd_sc_hd__clkbuf_2
X$15193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15195 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15199 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15200 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15201 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15202 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15205 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15206 VGND \$516 \$1289 \$1273 \$1288 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15207 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15208 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15209 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15211 VGND \$516 \$1275 \$1274 \$1290 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15213 VGND \$1261 \$1225 mgmt_gpio_out[2] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$15214 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15215 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15216 VPWR \$1291 VGND VPWR \$1393 \$1363 \$1261 \$1365 VGND
+ sky130_fd_sc_hd__o22a_1
X$15217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15222 VGND \$4473 \$3277 \$4493 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$15223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15224 VPWR \$4493 VGND VPWR \$4473 \$4508 \$1829 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$15225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15226 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15228 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15229 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15230 VPWR \$4441 VPWR VGND \$1979 \$3833 \$4474 VGND sky130_fd_sc_hd__or3_1
X$15231 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15233 VPWR \$4510 \$4351 VGND \$2511 VPWR \$4474 VGND sky130_fd_sc_hd__nor3_1
X$15234 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15235 VPWR \$4511 \$4265 VPWR \$1979 VGND \$3833 \$4210 VGND
+ sky130_fd_sc_hd__o211ai_1
X$15236 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15237 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15238 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15241 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15242 VGND \$4148 \$2214 \$4412 \$4512 \$4540 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$15243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15246 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15249 VPWR \$2215 \$4514 \$3693 VPWR VGND \$4513 \$4568 VGND
+ sky130_fd_sc_hd__or4_1
X$15250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15251 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15252 VPWR \$3637 \$4528 \$3157 VPWR VGND \$4527 \$4370 VGND
+ sky130_fd_sc_hd__or4_1
X$15253 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15254 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15255 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15256 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15257 VPWR \$4551 \$4516 \$4514 VPWR VGND \$4515 \$4529 VGND
+ sky130_fd_sc_hd__or4_1
X$15258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15260 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15261 VPWR \$4478 \$4309 \$4503 VPWR VGND \$4494 \$4486 VGND
+ sky130_fd_sc_hd__or4_1
X$15262 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15263 VPWR \$4487 VGND \$4504 \$4503 \$4432 VPWR \$3486 VGND
+ sky130_fd_sc_hd__nor4_1
X$15264 VPWR \$3776 \$4518 \$4486 VPWR VGND \$4517 \$4487 VGND
+ sky130_fd_sc_hd__or4_1
X$15265 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15266 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15267 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15268 VGND \$4447 \$4520 \$4519 \$4521 \$4157 \$4522 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$15269 VPWR \$4495 VPWR VGND \$3882 \$4486 \$4519 VGND sky130_fd_sc_hd__or3_2
X$15270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15273 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15274 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15275 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15276 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15277 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15278 VGND \$4374 \$4216 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$15279 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15280 VPWR VPWR VGND \$4255 \$4530 VGND sky130_fd_sc_hd__clkbuf_2
X$15281 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15282 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15283 VPWR VGND VPWR \$3251 \$4542 VGND sky130_fd_sc_hd__inv_2
X$15284 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15285 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15287 VPWR VGND \$4183 \$3711 \$4531 \$4532 \$4185 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15288 VPWR VGND VPWR \$4183 \$4185 VGND sky130_fd_sc_hd__inv_2
X$15289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15293 VPWR \$3999 \$4531 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15294 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15298 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15299 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15300 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15301 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15302 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15303 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15304 VGND \$4353 \$4534 \$4406 \$4533 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15305 VPWR VGND VPWR \$4405 \$4376 VGND sky130_fd_sc_hd__inv_2
X$15306 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15308 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15309 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15310 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15311 VGND \$4353 \$4489 \$4406 \$4488 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15312 VPWR \$3934 \$4534 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15313 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15314 VPWR VGND VPWR \$3963 \$4523 VGND sky130_fd_sc_hd__inv_2
X$15315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15316 VPWR VGND \$4407 \$3711 \$4489 \$4488 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15317 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15318 VGND \$4353 \$4496 \$4377 \$4524 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15319 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15320 VPWR VGND \$4407 \$1179 \$4496 \$4524 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15321 VPWR \$3746 \$4496 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15322 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15323 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15324 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15325 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15328 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15329 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15330 VPWR VGND VPWR \$4120 \$4497 VGND sky130_fd_sc_hd__inv_2
X$15331 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15333 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15335 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15336 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15337 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15339 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15340 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15342 VPWR VGND \$4407 \$354 \$4535 \$4536 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15344 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15347 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15348 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15349 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15350 VPWR \$4490 VGND VPWR \$3584 \$1625 \$4123 \$1466 VGND
+ sky130_fd_sc_hd__o22a_1
X$15351 VPWR VGND VPWR \$2629 \$4535 VGND sky130_fd_sc_hd__inv_2
X$15352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15353 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15354 VGND \$3727 \$4490 \$4087 \$2921 \$4239 \$4498 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15357 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15358 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15360 VGND \$3627 \$4525 \$4029 \$3019 \$2921 \$4279 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15364 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15365 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15366 VPWR \$4295 VGND VPWR \$4526 \$2919 \$4088 \$3019 VGND
+ sky130_fd_sc_hd__o22a_1
X$15367 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15370 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15372 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15374 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15375 VPWR VGND \$4357 \$1171 \$4497 \$4505 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15376 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15377 VGND \$2989 \$4497 \$4427 \$4505 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15380 VPWR \$4491 VGND \$2921 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$15381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15382 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15383 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15384 VPWR VGND \$4321 VPWR \$4491 VGND sky130_fd_sc_hd__clkbuf_4
X$15385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15388 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15389 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15390 VPWR \$4087 \$4500 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15391 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15392 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15393 VPWR VGND \$4303 \$411 \$4500 \$4506 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15394 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15395 VGND \$2989 \$4500 \$4165 \$4506 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15397 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15398 VGND \$2989 \$3297 \$4165 \$4537 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$15399 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15400 VPWR \$4537 VGND VPWR \$4547 \$4492 \$3297 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$15401 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15402 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15403 VPWR \$4472 VGND VPWR \$4775 \$4492 \$3738 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$15404 VGND \$2989 \$4167 \$4165 \$4502 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15405 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15407 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15408 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15412 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15413 VPWR VGND wb_dat_o[9] VPWR \$4438 VGND sky130_fd_sc_hd__buf_2
X$15414 VPWR VGND wb_dat_o[10] VPWR \$4473 VGND sky130_fd_sc_hd__buf_2
X$15415 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15418 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15420 VPWR \$4429 VPWR VGND \$1962 \$3833 \$4474 VGND sky130_fd_sc_hd__or3_1
X$15421 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15422 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15423 VPWR \$4429 \$4299 VPWR \$4439 VGND \$4440 \$3853 VGND
+ sky130_fd_sc_hd__o211ai_1
X$15424 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15425 VPWR \$4440 VGND VPWR \$4474 \$2511 \$4474 \$2552 VGND
+ sky130_fd_sc_hd__o22a_1
X$15426 VPWR \$4441 \$3805 VPWR \$4429 VGND VGND sky130_fd_sc_hd__and2_1
X$15427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15429 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15431 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15432 VPWR VPWR \$3856 VGND \$4475 \$4305 \$4419 \$4456 VGND
+ sky130_fd_sc_hd__a211o_1
X$15433 VGND \$4430 \$3918 \$4442 \$4443 \$3470 \$2001 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_2
X$15434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15436 VPWR VPWR \$2001 VGND \$4476 \$4411 \$4443 VGND sky130_fd_sc_hd__o21ai_1
X$15437 VGND \$4456 \$4431 \$4457 \$4305 \$4411 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$15438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15439 VPWR \$4431 VPWR VGND \$2742 \$1963 VGND sky130_fd_sc_hd__nand2_1
X$15440 VPWR VGND VPWR \$4457 \$4476 VGND sky130_fd_sc_hd__inv_2
X$15441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15442 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15443 VGND \$4457 \$4478 \$2257 \$4305 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$15444 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15445 VGND \$3859 \$4513 \$3709 \$4195 \$4444 \$4445 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_2
X$15446 VPWR VGND VPWR \$4420 \$4477 VGND sky130_fd_sc_hd__inv_2
X$15447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15448 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15449 VGND \$4468 \$4420 \$4457 \$2257 \$4458 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$15450 VGND \$4457 \$4458 \$4397 \$4420 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$15451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15453 VPWR \$4459 VGND \$4458 \$4398 VPWR VGND sky130_fd_sc_hd__or2_1
X$15454 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15455 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15457 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15458 VPWR \$4485 VPWR VGND \$4478 \$4468 \$4399 VGND sky130_fd_sc_hd__or3_1
X$15459 VPWR \$4486 VGND \$4432 \$4468 VPWR VGND sky130_fd_sc_hd__or2_1
X$15460 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15461 VPWR \$4433 VGND VPWR \$4446 VGND sky130_fd_sc_hd__clkbuf_1
X$15462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15463 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15465 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15466 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15467 VPWR VGND VPWR \$4421 \$4447 VGND sky130_fd_sc_hd__inv_2
X$15468 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15469 VPWR \$4434 VGND VPWR \$4516 VGND sky130_fd_sc_hd__clkbuf_1
X$15470 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15477 VGND \$2777 \$4383 \$4216 \$4435 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15480 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15481 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15483 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15484 VGND \$4353 \$4414 \$3921 \$4460 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15485 VPWR VGND \$4183 \$1179 \$4414 \$4460 \$4185 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15486 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15488 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15489 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15492 VGND \$4353 \$4448 \$3921 \$4461 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15493 VPWR VGND \$4270 \$3694 \$4448 \$4461 \$4272 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15495 VPWR \$3002 \$4448 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15497 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15499 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15500 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15502 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15504 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15506 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15509 VPWR \$3350 \$4489 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15511 VPWR VGND VPWR \$4407 \$4363 VGND sky130_fd_sc_hd__inv_2
X$15512 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15513 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15516 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15517 VGND \$4422 \$4449 \$4237 \$2358 \$2274 \$3721 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15519 VPWR \$4449 VGND VPWR \$3937 \$1954 \$3936 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15520 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15521 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15522 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15523 VGND \$4451 \$4450 \$3368 \$2358 \$2274 \$3527 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15524 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15525 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15526 VPWR \$4450 VGND VPWR \$3536 \$1954 \$4053 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15528 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15529 VGND \$4462 \$4451 \$3417 \$785 \$2220 \$3350 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15530 VGND \$3373 \$4499 \$3624 \$1561 \$3553 \$3514 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15532 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15533 VPWR \$4479 VGND VPWR \$3965 \$1954 \$3967 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15534 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15535 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15536 VGND \$4452 \$4479 \$4480 \$2358 \$2274 \$3476 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15538 VGND \$4292 \$4452 \$2600 \$785 \$2220 \$3746 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15539 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15540 VPWR \$4463 VGND VPWR \$2615 \$1954 \$2666 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15541 VGND \$4423 \$4463 \$2547 \$2358 \$2274 \$2691 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15542 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15543 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15545 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15546 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15548 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15549 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15550 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15551 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15552 VPWR \$4464 VGND VPWR \$2531 \$1954 \$4124 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15553 VPWR \$4469 VGND VPWR \$2854 \$1954 \$1821 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15554 VGND \$4425 \$4464 \$3944 \$2358 \$2274 \$3543 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15555 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15558 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15559 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15560 VGND \$4470 \$4469 \$4481 \$2358 \$2274 \$2863 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15561 VPWR \$4465 VGND VPWR \$2628 \$1954 \$3771 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$15562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15563 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15565 VGND \$4453 \$4465 \$4482 \$2358 \$2274 \$3518 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15566 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15567 VGND \$4454 \$4453 \$3782 \$785 \$2220 \$2629 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$15568 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15569 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15570 VGND \$4470 \$1949 \$785 \$2220 \$1855 \$2907 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$15571 VGND \$2989 \$4436 \$4164 \$4466 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15572 VPWR VGND VPWR \$3783 \$4436 VGND sky130_fd_sc_hd__inv_2
X$15573 VPWR VGND \$4357 \$354 \$4436 \$4466 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15575 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15576 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15579 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15580 VPWR \$4499 \$4483 VPWR \$4241 VGND \$2921 \$3924 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$15581 VPWR \$4241 \$4455 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15582 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15583 VGND \$2989 \$4455 \$4427 \$4467 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15584 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15585 VPWR VGND \$4303 \$386 \$4455 \$4467 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15588 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15589 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15592 VGND \$2989 \$3319 \$4165 \$4437 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$15593 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15594 VGND \$3952 \$4165 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$15595 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15597 VGND \$2989 \$3738 \$4165 \$4472 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15598 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15600 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15605 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15607 VPWR \$1367 VGND VPWR sram_ro_data[14] VGND sky130_fd_sc_hd__clkbuf_1
X$15608 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15611 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15613 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15614 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15615 VGND \$1431 \$1396 \$387 \$1409 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15616 VPWR \$1431 VGND VPWR \$1375 VGND sky130_fd_sc_hd__clkbuf_1
X$15617 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15618 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15619 VGND \$1432 \$1385 \$381 \$1410 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$15620 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15621 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15622 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15623 VPWR \$1441 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$15624 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15625 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15626 VPWR \$1432 VGND VPWR \$1441 VGND sky130_fd_sc_hd__clkbuf_1
X$15627 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15628 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15629 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15630 VPWR VGND \$1053 \$1442 \$1433 \$1397 \$1055 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15631 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15632 VPWR \$1416 VGND VPWR \$1377 VGND sky130_fd_sc_hd__clkbuf_1
X$15633 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15635 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15636 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15639 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15641 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15642 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15644 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15645 VGND \$1369 \$1387 \$2244 \$1379 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$15646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15647 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15648 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15649 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15651 VGND \$1018 \$1424 \$1378 \$482 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$15652 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15653 VPWR \$1424 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$15654 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15655 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15657 VPWR VGND VPWR \$1399 \$1417 VGND sky130_fd_sc_hd__inv_2
X$15658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15659 VPWR VGND \$1399 \$183 \$1418 \$1400 \$1417 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15660 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15661 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15662 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15663 VPWR VGND VPWR \$1419 \$1388 VGND sky130_fd_sc_hd__inv_2
X$15664 VGND \$1183 \$1385 \$1369 \$1452 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$15665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15666 VPWR \$1443 \$1418 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15668 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15670 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15671 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15672 VPWR \$1401 VGND VPWR \$1271 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15673 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15674 VPWR \$1444 VGND VPWR \$456 \$1034 VGND sky130_fd_sc_hd__or2_4
X$15675 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15676 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15677 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15678 VPWR \$1435 VGND VPWR \$1340 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15679 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15680 VPWR \$1318 \$1412 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15681 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15682 VGND \$1389 \$1257 \$1317 \$1412 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15683 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15684 VGND \$1389 \$1444 \$1317 \$1318 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15685 VGND \$1318 \$1425 \$1326 \$1389 \$1328 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15686 VGND \$1318 \$1435 \$1379 \$1389 \$1328 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15687 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15688 VGND \$1412 \$1434 \$1379 \$1389 \$1328 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15689 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15690 VGND \$1353 \$1445 \$1328 \$1412 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15691 VGND \$1353 \$1426 \$1328 \$1318 \$1326 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15692 VPWR VPWR VGND \$1446 \$463 VGND sky130_fd_sc_hd__clkbuf_2
X$15693 VGND \$1353 \$1454 \$1328 \$1412 \$1379 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15694 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15695 VPWR \$1435 VGND VPWR \$326 \$1034 VGND sky130_fd_sc_hd__or2_4
X$15696 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15697 VPWR \$1342 VGND VPWR \$923 \$1425 VGND sky130_fd_sc_hd__or2_4
X$15698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15699 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15700 VPWR \$1426 VGND VPWR \$1125 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15701 VPWR \$1034 VGND VPWR \$420 \$1425 VGND sky130_fd_sc_hd__or2_4
X$15702 VPWR \$1434 VGND VPWR \$520 \$1248 VGND sky130_fd_sc_hd__or2_4
X$15703 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15704 VPWR \$1264 VGND VPWR \$379 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15706 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15707 VPWR \$1329 VGND VPWR \$1089 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15708 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15709 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15710 VPWR \$1420 VGND VPWR \$1300 \$1342 VGND sky130_fd_sc_hd__or2_4
X$15711 VPWR \$1426 VGND VPWR \$320 \$1034 VGND sky130_fd_sc_hd__or2_4
X$15712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15714 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15716 VPWR \$1329 VGND VPWR \$188 \$1034 VGND sky130_fd_sc_hd__or2_4
X$15717 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15719 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15722 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15723 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15725 VPWR VGND VPWR \$1427 \$1358 VGND sky130_fd_sc_hd__inv_2
X$15726 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15728 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15729 VPWR \$1404 VGND \$1421 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$15730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15733 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15734 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15735 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15736 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15737 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15738 VGND \$1152 \$1422 \$1203 \$1436 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15739 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15740 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15741 VPWR VGND \$1303 \$354 \$1422 \$1436 \$1295 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15742 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15743 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15744 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15745 VPWR VGND \$1170 \$1179 \$1447 \$1437 \$1182 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15746 VGND \$297 \$264 \$188 \$1561 \$1423 \$1428 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$15747 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15748 VGND \$1152 \$1447 \$993 \$1437 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15749 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15750 VGND \$1152 \$1413 \$993 \$1391 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15752 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15753 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15754 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15756 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15757 VPWR \$1414 VGND VPWR \$1449 \$1448 VGND sky130_fd_sc_hd__or2_4
X$15758 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15759 VPWR \$1414 VGND VPWR \$1438 \$1374 VGND sky130_fd_sc_hd__or2_4
X$15760 VPWR VGND VPWR \$1448 \$1374 VGND sky130_fd_sc_hd__inv_2
X$15761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15762 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15763 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15764 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15766 VGND \$1406 \$464 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$15767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15769 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15770 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15773 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15775 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15776 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15778 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15779 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15780 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15781 VGND \$516 \$1450 \$1273 \$1439 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15782 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15784 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15786 VGND \$516 \$1430 \$1273 \$1429 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15787 VPWR VGND \$1311 \$542 \$1430 \$1429 \$1310 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15789 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15790 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15791 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15792 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15793 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15794 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15796 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15797 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15798 VPWR VGND wb_dat_o[16] VPWR \$4776 VGND sky130_fd_sc_hd__buf_2
X$15799 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15802 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15804 VPWR VGND \$3547 VPWR \$5214 VGND sky130_fd_sc_hd__clkbuf_4
X$15805 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15806 VGND \$2015 \$2336 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$15807 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15808 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15809 VPWR \$4211 VPWR VGND \$3833 \$3342 VGND sky130_fd_sc_hd__or2_2
X$15810 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15811 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15812 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15814 VPWR \$4602 VGND \$1897 \$4698 VPWR VGND sky130_fd_sc_hd__or2_1
X$15815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15817 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15819 VPWR \$4368 VGND \$4752 \$4214 VPWR VGND sky130_fd_sc_hd__or2_1
X$15820 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15821 VPWR \$4786 VGND \$4368 \$4061 VPWR VGND sky130_fd_sc_hd__or2_1
X$15822 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15825 VGND \$2257 \$4772 \$4663 \$4664 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$15826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15828 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15829 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15830 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15832 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15833 VPWR \$4778 VGND \$4777 \$4485 VPWR VGND sky130_fd_sc_hd__or2_1
X$15834 VPWR \$4310 VGND \$4752 \$4757 VPWR VGND sky130_fd_sc_hd__or2_1
X$15835 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15837 VPWR \$4787 VGND \$4778 \$4570 VPWR VGND sky130_fd_sc_hd__or2_1
X$15838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15839 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15840 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15841 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15842 VPWR \$4699 VGND \$4737 \$4758 VPWR VGND sky130_fd_sc_hd__or2_1
X$15843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15845 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15846 VPWR \$4572 VGND \$4727 \$4739 VPWR VGND sky130_fd_sc_hd__or2_1
X$15847 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15850 VPWR \$4773 VGND VPWR \$4789 VGND sky130_fd_sc_hd__clkbuf_1
X$15851 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15852 VGND \$3507 \$4779 \$4773 \$2082 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$15853 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15854 VPWR \$4741 VGND VPWR \$4759 VGND sky130_fd_sc_hd__clkbuf_1
X$15855 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15856 VPWR VGND VPWR \$4555 \$4530 VGND sky130_fd_sc_hd__inv_2
X$15857 VPWR VGND \$4555 \$293 \$4780 \$4812 \$4530 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15858 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15860 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15861 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15863 VPWR \$3814 \$4780 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15864 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15866 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15867 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15868 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15869 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15870 VPWR \$3642 \$4790 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$15871 VPWR VGND \$4760 \$3732 \$4703 \$4742 \$4717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15872 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15873 VGND \$4353 \$4761 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$15874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15875 VPWR \$1219 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$15876 VPWR \$4791 VGND \$1219 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$15877 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15880 VPWR VGND \$4781 \$1179 \$4704 \$4743 \$4782 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15881 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15882 VGND \$4353 \$4744 \$4406 \$4753 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15883 VPWR VGND \$4781 \$3694 \$4744 \$4753 \$4782 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15884 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15886 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15887 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15888 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15889 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15890 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15892 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15893 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15894 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15895 VPWR VPWR VGND \$4783 \$4374 VGND sky130_fd_sc_hd__clkbuf_2
X$15896 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15897 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15898 VGND \$4353 \$4745 \$4377 \$4762 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$15899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15900 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15901 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15902 VPWR VGND \$4707 \$1179 \$4745 \$4762 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15904 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15905 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15906 VGND \$4353 \$4754 \$4377 \$4763 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15908 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15909 VPWR VGND \$4707 \$3711 \$4754 \$4763 \$4706 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15910 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15911 VPWR VGND VPWR \$3923 \$4754 VGND sky130_fd_sc_hd__inv_2
X$15912 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15915 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15916 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15917 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15918 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15919 VGND \$4353 \$4764 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$15920 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15921 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15922 VPWR VGND \$4681 \$542 \$4226 \$4755 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15924 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15925 VGND \$4353 \$4226 \$4424 \$4755 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$15926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15928 VGND \$4353 \$4747 \$4424 \$4748 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15929 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15930 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15931 VPWR VGND \$4681 \$411 \$4784 \$4793 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15932 VPWR VGND VPWR \$1893 \$4784 VGND sky130_fd_sc_hd__inv_2
X$15933 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15934 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15935 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15936 VPWR VGND \$4681 \$184 \$4756 \$4766 \$4682 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15937 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15938 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15939 VGND \$4353 \$4756 \$4765 \$4766 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15940 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15941 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15942 VPWR \$4794 VGND \$2918 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$15943 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15944 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15945 VPWR \$4795 VGND \$2751 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$15946 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$15947 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15949 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15950 VPWR \$4767 VGND \$3121 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$15951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15953 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15954 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15955 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15956 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15960 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15963 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15964 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15965 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15966 VPWR VGND \$4750 \$1677 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$15967 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15968 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15969 VGND \$2989 \$4751 \$4165 \$4768 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15970 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15971 VPWR \$4768 VGND VPWR \$4769 \$4492 \$4751 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$15972 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15973 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15976 VPWR VGND \$4650 \$1179 \$4785 \$4770 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$15977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15978 VGND \$4775 \$1179 \$4785 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$15979 VGND \$2989 \$4785 \$4165 \$4770 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$15980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15981 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$15983 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15984 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15985 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15986 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$15987 VGND \$3279 \$3277 \$3278 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$15988 VGND spi_sck \$3247 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$15989 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15991 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$15992 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$15993 VGND \$3248 \$3255 \$3231 \$2939 \$3140 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$15994 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$15996 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15997 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$15998 VPWR \$3257 VPWR VGND \$3256 \$3173 \$2388 VGND sky130_fd_sc_hd__or3b_1
X$15999 VPWR \$3258 VGND \$3115 \$3173 VPWR VGND sky130_fd_sc_hd__or2_1
X$16000 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16001 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16002 VPWR \$3256 \$3268 \$3267 VPWR VGND \$3100 \$2925 VGND
+ sky130_fd_sc_hd__or4_1
X$16003 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16004 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16005 VPWR \$3232 VGND \$2817 \$3268 VPWR VGND sky130_fd_sc_hd__or2_1
X$16006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16007 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16008 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16009 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16010 VPWR VGND \$2514 VPWR \$3249 VGND sky130_fd_sc_hd__clkbuf_4
X$16011 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16012 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16013 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16014 VGND \$3175 \$3260 \$3259 \$2643 \$2639 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$16015 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16016 VPWR VGND \$2488 VPWR \$3280 VGND sky130_fd_sc_hd__clkbuf_4
X$16017 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16018 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16019 VPWR \$2741 \$3269 \$2488 \$3141 VGND \$2996 VPWR VGND
+ sky130_fd_sc_hd__o22ai_1
X$16020 VPWR \$3281 VGND \$3269 \$3233 VPWR VGND sky130_fd_sc_hd__or2_1
X$16021 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16022 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16023 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16024 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16025 VPWR \$3261 VGND \$3176 \$3250 VPWR VGND sky130_fd_sc_hd__or2_1
X$16026 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16027 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16028 VPWR \$3250 VGND \$2472 VPWR \$2949 VGND sky130_fd_sc_hd__nor2_1
X$16029 VPWR \$3282 VGND \$3250 \$3119 VPWR VGND sky130_fd_sc_hd__or2_1
X$16030 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16031 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16032 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16033 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16034 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16035 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16036 VGND \$2777 \$3270 \$2556 \$3283 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16037 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16038 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16039 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16040 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16041 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16042 VPWR VGND \$3284 \$183 \$3285 \$3306 \$3304 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16046 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16047 VPWR \$2936 \$3285 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16050 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16051 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16052 VPWR VPWR VGND \$3286 \$2954 VGND sky130_fd_sc_hd__clkbuf_2
X$16053 VPWR \$3144 \$3158 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16057 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16058 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16061 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16062 VPWR \$1570 VGND VPWR \$3271 \$1435 VGND sky130_fd_sc_hd__or2_4
X$16063 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16064 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16065 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16066 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16067 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16068 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16069 VPWR \$3220 VGND VPWR \$2999 \$3106 \$3002 \$3271 VGND
+ sky130_fd_sc_hd__o22a_1
X$16070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16071 VGND \$3072 \$3234 \$3262 \$2830 \$2651 \$3251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16072 VPWR \$3219 VGND VPWR \$3251 \$2254 \$2971 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$16073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16074 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16076 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16077 VPWR \$3160 VGND \$2007 \$3262 VPWR VGND sky130_fd_sc_hd__or2_1
X$16078 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16079 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16081 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16082 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16083 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16084 VPWR wb_clk_i VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16086 VGND wb_clk_i \$3133 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$16087 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16088 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16090 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16091 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16092 VPWR VGND VPWR \$3291 \$3290 \$3145 \$3288 \$3289 VGND
+ sky130_fd_sc_hd__and4_1
X$16093 VPWR \$3221 VGND VPWR \$3131 \$2734 \$3122 \$2789 VGND
+ sky130_fd_sc_hd__o22a_1
X$16094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16096 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16097 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16098 VPWR \$3264 VGND VPWR \$3263 \$1956 \$2191 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$16099 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16100 VGND \$3272 \$2725 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$16101 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16102 VGND \$3237 \$3329 \$2900 \$2830 \$2651 \$2502 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16103 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16104 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16105 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16106 VPWR \$3186 VGND VPWR \$2163 \$1967 \$3265 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$16107 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16108 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16109 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16111 VGND \$3252 \$3253 \$3239 \$3044 VPWR \$1127 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$16112 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16113 VGND \$4317 \$3240 \$2252 \$2047 \$2048 \$3292 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16115 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16117 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16118 VPWR \$3167 VGND VPWR \$1720 \$1300 \$3254 \$2162 VGND
+ sky130_fd_sc_hd__o22a_1
X$16119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16121 VPWR \$3273 VGND VPWR \$731 \$2045 \$2813 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$16122 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16123 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16125 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16126 VGND \$3274 \$1880 \$2005 \$3336 \$3293 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$16127 VPWR \$3226 VGND VPWR \$3254 \$1967 \$3465 \$1939 VGND
+ sky130_fd_sc_hd__o22a_1
X$16128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16130 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16131 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16132 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16133 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16134 VPWR VGND VPWR \$3225 \$3210 \$3656 \$3243 \$3211 VGND
+ sky130_fd_sc_hd__and4_1
X$16135 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16136 VPWR \$3275 VGND VPWR \$3294 \$1956 \$2053 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$16137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16138 VPWR \$3266 VGND VPWR \$3111 \$1956 \$2307 \$1957 VGND
+ sky130_fd_sc_hd__o22a_1
X$16139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16142 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16144 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16145 VPWR VGND VPWR \$3294 \$3150 VGND sky130_fd_sc_hd__inv_2
X$16146 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16149 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16150 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16151 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16153 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16154 VPWR \$3328 \$3244 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16155 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16157 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16158 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16159 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16161 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16162 VPWR VGND \$3169 \$354 \$3296 \$3295 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16163 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16166 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16167 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16169 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16170 VPWR VGND VPWR \$3169 \$3171 VGND sky130_fd_sc_hd__inv_2
X$16171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16172 VGND \$3276 \$1333 \$3297 \$741 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16173 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16174 VGND \$3276 \$2829 mgmt_gpio_out[8] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$16175 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16176 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16177 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16179 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16181 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16182 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16183 VPWR VGND sram_ro_addr[7] VPWR \$484 VGND sky130_fd_sc_hd__buf_2
X$16184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16189 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16190 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16192 VPWR \$491 \$513 VPWR \$462 VGND \$481 VGND sky130_fd_sc_hd__o21ba_1
X$16193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16197 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16199 VGND \$537 \$440 \$381 \$536 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16200 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16201 VPWR \$537 VGND VPWR \$544 VGND sky130_fd_sc_hd__clkbuf_1
X$16202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16204 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16206 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16207 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16208 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16210 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16212 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16213 VGND \$655 \$182 \$237 \$505 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$16214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16216 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16218 VPWR VGND VPWR \$524 \$182 VGND sky130_fd_sc_hd__inv_2
X$16219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16220 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16222 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16223 VPWR VGND \$525 VPWR \$546 VGND sky130_fd_sc_hd__buf_2
X$16224 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16225 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16226 VPWR \$546 VGND \$1103 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$16227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16228 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16231 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16233 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16234 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16236 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16237 VPWR VGND \$514 \$294 \$486 \$494 \$515 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16238 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16239 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16240 VGND \$206 \$516 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$16241 VPWR VGND VPWR \$514 \$515 VGND sky130_fd_sc_hd__inv_2
X$16242 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16243 VPWR VGND \$514 \$183 \$547 \$559 \$515 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16244 VPWR VGND \$486 \$495 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$16245 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16246 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16247 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16248 VGND \$463 \$196 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$16249 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16250 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16251 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16252 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16253 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16254 VGND \$517 \$507 \$320 \$457 \$520 \$572 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_4
X$16255 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16256 VGND \$516 \$528 \$198 \$548 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16257 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16258 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16259 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16260 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16261 VGND \$516 \$569 \$198 \$549 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16264 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16265 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16267 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16268 VPWR \$497 VGND VPWR \$495 \$1266 \$190 \$188 VGND
+ sky130_fd_sc_hd__o22a_1
X$16269 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16271 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16273 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16274 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16275 VGND \$529 \$509 \$326 \$686 \$485 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$16276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16277 VGND \$206 \$518 \$435 \$530 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16280 VPWR VGND \$417 \$293 \$518 \$530 \$434 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16282 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16285 VPWR \$512 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16286 VPWR \$512 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16287 VGND \$421 \$348 \$512 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16288 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16289 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16290 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16291 VPWR \$512 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16293 VGND \$426 \$406 \$487 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16294 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16295 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16297 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16298 VPWR \$526 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16299 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16300 VGND \$511 \$406 \$526 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16301 VPWR \$519 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16302 VGND \$330 \$399 \$519 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16303 VGND \$502 \$399 \$540 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16304 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16306 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16307 VPWR \$540 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16308 VPWR VGND \$417 \$184 \$550 \$561 \$434 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16309 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16310 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16311 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16312 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16313 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16314 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16315 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16316 VGND \$501 \$289 \$459 \$532 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$16317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16318 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16321 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16322 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16323 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16325 VGND \$468 \$289 \$480 \$510 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$16326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16329 VGND \$206 \$562 \$541 \$551 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16330 VPWR \$521 VGND \$520 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$16331 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16332 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16334 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16335 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16336 VPWR VGND \$292 VPWR \$521 VGND sky130_fd_sc_hd__buf_2
X$16337 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16338 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16339 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16340 VGND \$294 \$534 \$533 \$291 \$292 VPWR VPWR VGND
+ sky130_fd_sc_hd__a22o_2
X$16341 VGND \$206 \$534 \$254 \$533 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$16342 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16343 VPWR VGND \$291 \$542 \$552 \$543 \$292 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16344 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16345 VGND \$206 \$552 \$254 \$543 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$16346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16347 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16350 VPWR VGND \$211 \$553 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$16351 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16352 VGND mgmt_gpio_in[0] \$2550 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$16353 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16355 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16356 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16357 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16359 VPWR \$3278 VGND VPWR \$3279 \$3531 \$907 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$16360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16361 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16362 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16365 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16367 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16368 VPWR VGND \$3501 \$2944 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$16369 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16370 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16373 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16374 VPWR VGND VPWR \$3548 \$3487 VGND sky130_fd_sc_hd__inv_2
X$16375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16376 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16377 VPWR \$2663 \$3550 \$3549 VPWR VGND \$3117 \$2444 VGND
+ sky130_fd_sc_hd__or4_1
X$16378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16379 VGND \$3493 \$3499 \$3573 \$3521 \$3780 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$16380 VPWR \$3506 VGND VPWR \$3503 VGND sky130_fd_sc_hd__clkbuf_1
X$16381 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16382 VPWR VGND VPWR \$3521 \$3550 VGND sky130_fd_sc_hd__inv_2
X$16383 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16387 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16388 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16393 VPWR \$1831 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16394 VGND \$3532 \$1831 \$2330 \$2219 \$3551 \$2105 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$16395 VPWR \$3552 VGND VPWR \$3180 \$1954 \$3508 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$16396 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16397 VPWR \$3522 VGND VPWR \$3144 \$2456 \$3349 \$2416 VGND
+ sky130_fd_sc_hd__o22a_1
X$16398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16399 VGND \$3459 \$3533 \$712 \$785 \$2220 \$3144 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16401 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16402 VGND \$3495 \$3510 \$712 \$2369 \$2357 \$3348 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16403 VGND \$3511 \$3565 \$3508 \$2750 \$2541 \$646 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16405 VPWR \$3523 VGND \$3553 \$2664 VPWR VGND sky130_fd_sc_hd__or2_1
X$16406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16407 VPWR \$2550 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16408 VPWR VGND VPWR \$3554 \$2550 VGND sky130_fd_sc_hd__inv_2
X$16409 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16410 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16411 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16412 VGND \$3555 \$3534 \$3263 \$2325 \$3556 \$2611 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16413 VGND \$3461 \$3535 \$1265 \$1271 \$2375 \$3536 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16414 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16415 VPWR \$1646 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16416 VGND \$3372 \$1646 \$3537 \$2734 \$1676 \$3538 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16417 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16418 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16420 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16421 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16422 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16423 VGND \$3539 \$3488 \$2994 \$2785 \$1839 \$3524 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16425 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16426 VPWR \$3526 VGND VPWR \$3540 \$2665 \$2397 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$16427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16428 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16429 VGND \$3253 \$3525 \$3527 \$2544 \$2545 \$3351 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16431 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16432 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16433 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16434 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16436 VPWR \$3336 VGND VPWR \$3541 \$2670 \$1702 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$16437 VGND \$3316 \$3542 \$3543 \$2544 \$2545 \$3496 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16439 VPWR \$3528 VGND VPWR \$3544 \$1966 \$3405 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$16440 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16441 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16442 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16443 VGND \$3545 \$3528 \$2605 \$2043 \$1914 \$3354 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16444 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16445 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16446 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16447 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16448 VPWR \$3520 VGND \$1839 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$16449 VPWR \$2587 \$3546 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16450 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16451 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16452 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16454 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16455 VGND \$1363 \$345 \$3568 \$927 \$4239 VPWR VPWR VGND
+ sky130_fd_sc_hd__a211o_4
X$16456 VPWR VGND \$3169 \$1171 \$3529 \$3557 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16457 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16458 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16459 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16460 VPWR VGND \$3169 \$1179 \$3530 \$3558 \$3171 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16461 VPWR \$3524 \$3530 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16462 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16463 VGND \$3739 mgmt_gpio_out[9] \$2791 VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_2
X$16464 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16465 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16466 VGND \$3592 \$3277 \$3591 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$16467 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16468 VGND \$3593 \$3571 \$3570 \$3139 VPWR VPWR \$2911 VGND
+ sky130_fd_sc_hd__or4b_1
X$16469 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16470 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16471 VPWR \$2363 \$3503 \$2169 VPWR VGND \$3571 \$3594 VGND
+ sky130_fd_sc_hd__or4_1
X$16472 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16473 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16474 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16475 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16477 VPWR \$3595 VGND \$2390 \$3596 VPWR VGND sky130_fd_sc_hd__or2_1
X$16478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16481 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16482 VPWR \$3779 VGND \$2966 \$3548 VPWR VGND sky130_fd_sc_hd__or2_1
X$16483 VPWR \$3549 VPWR VGND \$3572 \$3560 \$3302 VGND sky130_fd_sc_hd__or3_1
X$16484 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16485 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16486 VPWR VPWR \$3550 VGND \$3498 \$3561 \$3573 VGND sky130_fd_sc_hd__o21ai_1
X$16487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16488 VGND \$1741 \$3597 \$3598 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$16489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16492 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16495 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16496 VPWR \$2983 \$3574 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16497 VPWR \$1490 VGND VPWR \$3562 \$1059 VGND sky130_fd_sc_hd__or2_4
X$16498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16499 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16500 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16501 VPWR \$3532 VGND VPWR \$3564 \$2229 \$3563 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$16502 VPWR VGND VPWR \$3563 \$3641 VGND sky130_fd_sc_hd__inv_2
X$16503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16504 VGND \$3533 \$3552 \$3642 \$2358 \$2274 \$3509 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16506 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16507 VPWR \$1490 VGND VPWR \$3553 \$1434 VGND sky130_fd_sc_hd__or2_4
X$16508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16509 VPWR \$3565 VGND VPWR \$868 \$2559 \$3575 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$16510 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16511 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16512 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16513 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16514 VGND \$3149 \$3035 \$3553 \$3562 \$3251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$16515 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16516 VGND \$3599 \$3576 \$3554 \$927 \$2734 \$2477 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16517 VGND \$3600 \$3523 \$3328 \$1879 \$3106 \$2072 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16518 VGND \$899 \$3577 \$3578 VPWR \$1523 VPWR VGND sky130_fd_sc_hd__nand3_4
X$16519 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16520 VPWR \$3579 VGND VPWR \$3601 \$1966 \$2784 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$16521 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16522 VGND \$3580 \$3579 \$2841 \$2043 \$1914 \$3328 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16523 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16524 VPWR \$3566 VGND VPWR \$3581 \$2670 \$1071 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$16525 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16526 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16527 VGND \$3622 \$3567 \$1820 \$1890 \$1561 \$3601 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16530 VPWR \$3525 VGND VPWR \$3538 \$2665 \$4107 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$16531 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16532 VGND \$3603 \$3602 \$2400 \$2043 \$1914 \$3378 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16533 VGND \$3604 \$3582 \$3351 \$2043 \$1914 \$1927 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16535 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16536 VPWR VGND VPWR \$3606 \$3583 \$3449 \$3605 \$2431 VGND
+ sky130_fd_sc_hd__and4_1
X$16537 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16538 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16539 VPWR \$3542 VGND VPWR \$1893 \$2665 \$3584 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$16540 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16541 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16542 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16543 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16544 VGND \$3607 \$3585 \$2756 \$927 \$1676 \$3586 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16545 VPWR \$3517 VGND VPWR \$3586 \$2665 \$3587 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$16546 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16549 VGND \$3608 \$3657 \$3467 \$2043 \$1914 \$3112 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16550 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16551 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16553 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16554 VPWR \$3567 \$3588 VPWR \$269 VGND \$1562 \$3609 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$16555 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16556 VGND \$2989 \$3546 \$3425 \$3610 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16559 VPWR VGND \$3589 \$2791 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$16560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16561 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16562 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16563 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16564 VGND \$3568 \$3611 \$1335 \$1083 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16566 VGND \$2989 \$3529 \$3425 \$3557 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16567 VGND \$2989 \$3530 \$3590 \$3558 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16568 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16569 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16570 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16571 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16573 VGND \$3740 \$3277 \$3757 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$16574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16575 VPWR \$3757 VGND VPWR \$3740 \$3531 \$1829 \$3547 VGND
+ sky130_fd_sc_hd__o22a_1
X$16576 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16577 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16578 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16579 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16580 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16581 VGND \$2320 \$3854 \$3357 \$3470 \$2571 \$3742 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_4
X$16582 VGND \$3758 \$2336 \$1998 \$3057 \$3690 \$3741 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$16583 VPWR \$3689 VGND \$3742 VPWR \$2741 VGND sky130_fd_sc_hd__nor2_1
X$16584 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16586 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16588 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16589 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16591 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16592 VPWR \$2940 \$3807 \$3199 VPWR VGND \$3759 \$3806 VGND
+ sky130_fd_sc_hd__or4_1
X$16593 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16594 VPWR \$3175 \$3775 VGND \$2940 VPWR \$3776 \$3787 VGND
+ sky130_fd_sc_hd__or4_2
X$16595 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16598 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16599 VPWR \$3473 \$3778 \$3777 VPWR VGND \$3787 \$3260 VGND
+ sky130_fd_sc_hd__or4_1
X$16600 VPWR \$3808 VPWR VGND \$3281 \$3779 \$3788 VGND sky130_fd_sc_hd__or3_1
X$16601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16603 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16604 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16605 VPWR \$3809 VPWR VGND \$3789 \$3343 \$2978 VGND sky130_fd_sc_hd__or3b_1
X$16606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16609 VGND \$3780 \$3807 \$3790 \$3791 \$3792 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$16610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16611 VPWR VGND VPWR \$3791 \$3778 VGND sky130_fd_sc_hd__inv_2
X$16612 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16613 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16615 VPWR VGND VPWR \$3810 \$3793 VGND sky130_fd_sc_hd__inv_2
X$16616 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16617 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16619 VPWR VGND \$3667 \$3732 \$3812 \$3811 \$3669 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16620 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16621 VGND \$2777 \$3684 \$3413 \$3731 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16622 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16623 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16624 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16625 VGND \$3813 \$3413 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$16626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16627 VGND \$856 \$3743 \$3413 \$3760 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16629 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16630 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16631 VPWR VGND \$3435 \$3732 \$3743 \$3760 \$3458 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16632 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16633 VGND \$856 \$3761 \$3413 \$3733 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16634 VPWR VGND \$3435 \$293 \$3761 \$3733 \$3458 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16635 VPWR VGND VPWR \$3713 \$3743 VGND sky130_fd_sc_hd__inv_2
X$16636 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16637 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16638 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16639 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16640 VPWR VGND VPWR \$3719 \$3761 VGND sky130_fd_sc_hd__inv_2
X$16641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16642 VPWR \$3744 VGND VPWR \$3840 \$2229 \$3713 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$16643 VGND \$2801 \$3744 \$2644 \$2330 \$2219 \$3864 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16645 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16646 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16647 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16648 VPWR \$1570 VGND VPWR \$3556 \$1425 VGND sky130_fd_sc_hd__or2_4
X$16649 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16650 VPWR \$3762 VGND VPWR \$3712 \$2927 \$818 \$2616 VGND
+ sky130_fd_sc_hd__o22a_1
X$16651 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16652 VGND \$2542 \$3762 \$3734 \$2830 \$2651 \$3814 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16653 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16654 VPWR \$3763 VGND VPWR \$2296 \$2366 \$3734 \$3204 VGND
+ sky130_fd_sc_hd__o22a_1
X$16655 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16656 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16657 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16658 VPWR \$3745 VGND \$2007 \$3704 VPWR VGND sky130_fd_sc_hd__or2_1
X$16659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16660 VGND \$3745 \$2664 \$2116 \$1536 \$1837 \$2138 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$16661 VPWR \$1060 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16662 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16663 VPWR \$3311 VGND VPWR \$3719 \$3143 \$3746 \$1819 VGND
+ sky130_fd_sc_hd__o22a_1
X$16664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16665 VPWR \$1019 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16666 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16668 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16669 VPWR \$2671 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16670 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16671 VPWR \$3815 VGND VPWR \$2671 \$2785 \$3216 \$3703 VGND
+ sky130_fd_sc_hd__o22a_1
X$16672 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16673 VGND \$3764 \$3720 \$3061 \$2785 \$3703 \$3564 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16674 VGND \$3088 \$3815 \$2866 \$3765 \$3556 \$3017 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16675 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16676 VPWR \$1570 VGND VPWR \$3765 \$1426 VGND sky130_fd_sc_hd__or2_4
X$16677 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16678 VPWR \$3747 VGND \$2007 \$3162 VPWR VGND sky130_fd_sc_hd__or2_1
X$16679 VGND \$3817 \$3074 \$3794 \$1715 \$1754 \$1242 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16680 VGND \$3766 \$3747 \$1730 \$2116 \$1536 \$1071 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16681 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16682 VPWR VGND VPWR \$3818 \$3817 \$3766 \$3580 \$3795 VGND
+ sky130_fd_sc_hd__and4_1
X$16683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16684 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16685 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16686 VGND \$3767 \$3763 \$3292 \$2581 \$1558 \$1239 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16687 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16688 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16689 VGND \$3767 \$3820 \$3797 \$3819 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$16690 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16691 VPWR VGND VPWR \$3821 \$3816 \$3539 \$2805 \$3798 VGND
+ sky130_fd_sc_hd__and4_1
X$16692 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16693 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16694 VPWR \$3821 \$3781 \$3820 VGND VPWR \$1703 VGND sky130_fd_sc_hd__and3_2
X$16695 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16697 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16698 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16699 VPWR \$3822 VGND VPWR \$3524 \$2254 \$3796 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$16700 VPWR VPWR VGND \$2725 \$3769 VGND sky130_fd_sc_hd__clkbuf_2
X$16701 VGND \$3823 \$2251 \$3748 \$2921 \$1879 \$3378 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16703 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16704 VGND \$3749 \$3822 \$1616 \$2809 \$3218 \$3748 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16705 VPWR VGND VPWR \$3770 \$3706 \$3725 \$3603 \$3749 VGND
+ sky130_fd_sc_hd__and4_1
X$16706 VGND \$3725 \$3750 \$3540 \$2116 \$1536 \$1644 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16707 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16708 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16709 VPWR \$3401 VGND VPWR \$3796 \$2670 \$1644 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$16710 VPWR \$1469 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16711 VGND \$3583 \$1469 \$3782 \$1466 \$1845 \$3771 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16712 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16713 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16714 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16715 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16716 VGND \$1883 \$3751 \$3728 \$3847 VPWR \$1769 VPWR VGND
+ sky130_fd_sc_hd__nand4_4
X$16717 VGND \$3824 \$3799 \$2813 \$2785 \$3121 \$3825 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16718 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16720 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16721 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16722 VPWR \$3585 VGND VPWR \$3783 \$2031 \$3752 \$2789 VGND
+ sky130_fd_sc_hd__o22a_1
X$16723 VGND \$3753 \$3686 \$3752 \$1715 \$1754 \$1390 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16724 VGND \$3827 \$3708 \$3782 \$2369 \$2357 \$3629 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16726 VPWR \$3826 VGND VPWR \$3783 \$2559 \$2430 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$16727 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16728 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16729 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16730 VPWR \$3800 VGND \$2007 \$3828 VPWR VGND sky130_fd_sc_hd__or2_1
X$16731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16732 VGND \$3754 \$3800 \$3586 \$2116 \$1536 \$2630 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16733 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16734 VPWR VGND VPWR \$3736 \$3753 \$3754 \$3545 \$3735 VGND
+ sky130_fd_sc_hd__and4_1
X$16735 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16736 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16737 VPWR \$3772 VGND VPWR \$3338 \$2254 \$3450 \$2590 VGND
+ sky130_fd_sc_hd__o22a_1
X$16738 VPWR \$3801 VGND VPWR \$3450 \$3765 \$3628 \$2581 VGND
+ sky130_fd_sc_hd__o22a_1
X$16739 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16740 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16741 VGND \$3784 \$3801 \$3518 \$2751 \$3121 \$3828 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$16742 VPWR \$3005 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16743 VPWR \$3844 \$3755 VPWR \$3005 VGND \$2180 \$3609 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$16744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16745 VPWR VGND \$3630 \$354 \$3802 \$3829 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16748 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16749 VPWR VGND VPWR \$3222 \$3737 VGND sky130_fd_sc_hd__inv_2
X$16750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16751 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16752 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16753 VGND \$2989 \$3737 \$3425 \$3773 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16754 VPWR VGND \$3630 \$386 \$3737 \$3773 \$3631 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16756 VPWR VGND VPWR \$2430 \$3730 VGND sky130_fd_sc_hd__inv_2
X$16757 VGND \$2989 \$3730 \$3425 \$3729 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16758 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16759 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16760 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16761 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16762 VPWR VGND VPWR \$3716 \$3717 VGND sky130_fd_sc_hd__inv_2
X$16763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16764 VPWR VGND \$3716 \$1594 \$3697 \$3718 \$3717 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16765 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16766 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16767 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16768 VPWR VGND VPWR \$3450 \$3803 VGND sky130_fd_sc_hd__inv_2
X$16769 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16770 VGND \$2989 \$3803 \$3590 \$3785 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16771 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16773 VPWR \$3796 \$3756 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16774 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16775 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16776 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16777 VPWR \$3738 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16778 VPWR \$3786 VGND VPWR \$3804 VGND sky130_fd_sc_hd__clkbuf_1
X$16779 VGND \$3739 \$4106 \$3738 \$482 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16780 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16781 VPWR \$3804 VGND VPWR \$2846 VGND sky130_fd_sc_hd__clkbuf_1
X$16782 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16783 VPWR VGND mgmt_gpio_oeb[10] VPWR \$3786 VGND sky130_fd_sc_hd__buf_2
X$16784 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16785 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16786 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16790 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16791 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16792 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16793 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16794 VPWR \$1091 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$16795 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16796 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16797 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16798 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16799 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16800 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16801 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16802 VPWR \$5493 VPWR VGND \$5647 \$5632 \$5646 VGND sky130_fd_sc_hd__or3b_1
X$16803 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16804 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16805 VGND \$5646 \$4916 \$4891 \$5606 \$5619 VPWR VPWR VGND
+ sky130_fd_sc_hd__a2bb2o_1
X$16806 VPWR VGND VPWR \$5632 \$5449 VGND sky130_fd_sc_hd__inv_2
X$16807 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16808 VPWR \$5147 VPWR VGND \$5449 \$4880 \$5633 VGND sky130_fd_sc_hd__or3_2
X$16809 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16810 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16811 VPWR \$5607 VGND VPWR \$4880 \$5633 \$4853 \$5619 VGND
+ sky130_fd_sc_hd__o22a_1
X$16812 VPWR VGND \$5509 VPWR \$4863 \$5628 \$5619 VGND sky130_fd_sc_hd__a21oi_1
X$16813 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16814 VPWR \$5607 VGND VPWR \$4078 \$5628 VGND sky130_fd_sc_hd__or2_4
X$16815 VPWR VGND VPWR \$5619 \$5633 VGND sky130_fd_sc_hd__inv_2
X$16816 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16817 VPWR VGND VPWR \$5597 \$5628 VGND sky130_fd_sc_hd__inv_2
X$16818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16819 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16820 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16821 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16822 VPWR VGND VPWR \$5618 \$5458 VGND sky130_fd_sc_hd__inv_2
X$16823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16825 VGND \$5608 \$5609 \$4106 \$5634 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16826 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16828 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16829 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16830 VPWR VGND \$5504 \$780 \$5609 \$5634 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16832 VGND \$4774 \$5609 \$1369 \$5648 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$16833 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16835 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16836 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16837 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16838 VGND \$3694 \$5496 \$1369 \$5686 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$16839 VGND \$5611 \$5575 \$4106 \$5639 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16841 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16842 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16843 VGND \$184 \$5575 \$1369 \$5649 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$16844 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16845 VGND \$411 \$5485 \$1369 \$5651 VPWR VPWR VGND sky130_fd_sc_hd__mux2_8
X$16846 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16847 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16849 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16850 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16851 VPWR VGND \$5620 VPWR \$5613 \$5592 \$5339 VGND sky130_fd_sc_hd__a21oi_1
X$16852 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16853 VPWR VPWR \$5567 VGND \$5586 \$5495 \$5621 \$5622 VGND
+ sky130_fd_sc_hd__a211o_1
X$16854 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16855 VGND \$5613 \$5621 \$5614 \$5423 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$16856 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16857 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16858 VGND \$5620 \$5622 \$5613 \$5079 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$16859 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16860 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16861 VPWR VGND VPWR \$5192 \$4803 VGND sky130_fd_sc_hd__inv_2
X$16862 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16863 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16864 VGND \$3732 \$1594 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$16865 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16866 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16867 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16870 VGND \$4023 \$1171 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$16871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16872 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16873 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16875 VGND \$2777 \$5623 \$5408 \$5635 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16876 VPWR VGND \$5388 \$4774 \$5623 \$5635 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16877 VGND \$4374 \$5408 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$16878 VPWR VGND VPWR \$5623 \$1612 VGND sky130_fd_sc_hd__inv_4
X$16879 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16880 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16882 VGND \$2777 \$5624 \$5408 \$5640 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16884 VPWR VGND \$5229 \$4774 \$5624 \$5640 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16886 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16887 VGND \$2777 \$5625 \$4994 \$5641 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16888 VPWR VGND \$5525 \$4774 \$5625 \$5641 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16889 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16890 VPWR VGND VPWR \$5625 \$2397 VGND sky130_fd_sc_hd__inv_4
X$16891 VPWR \$910 \$5624 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$16892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16893 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16894 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16895 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16896 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16897 VGND \$2777 \$5602 \$5367 \$5615 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$16898 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16901 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16902 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16903 VPWR VGND \$5562 \$1594 \$5601 \$5636 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16904 VGND \$4761 \$5601 \$5367 \$5636 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16906 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16907 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16908 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16909 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16910 VPWR VGND VPWR \$3584 \$5629 VGND sky130_fd_sc_hd__inv_2
X$16911 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16912 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16913 VGND \$4761 \$5626 \$5369 \$5642 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16914 VPWR VGND \$5562 \$411 \$5626 \$5642 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16915 VPWR VGND \$5626 \$2481 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$16916 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16917 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16920 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16921 VGND \$4761 \$5630 \$5272 \$5643 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16923 VPWR VGND \$5627 \$4774 \$5630 \$5643 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$16924 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16925 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16926 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16927 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16928 VGND \$4761 \$5664 \$5334 \$5644 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16929 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16930 VGND \$5595 \$5940 \$3609 \$2356 \$3611 VPWR VPWR VGND
+ sky130_fd_sc_hd__a22oi_4
X$16931 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16932 VGND \$5941 \$5616 \$3611 \$4320 \$3609 VPWR VPWR VGND
+ sky130_fd_sc_hd__a22oi_4
X$16933 VPWR VGND VPWR \$5627 \$5589 VGND sky130_fd_sc_hd__inv_2
X$16934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16935 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16937 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16938 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16939 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16940 VGND \$4764 \$5658 \$5298 \$5645 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$16941 VGND \$5579 \$1221 mgmt_gpio_out[31] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$16942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16943 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16944 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16945 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16946 VPWR \$5650 VGND VPWR \$5637 \$4724 \$5652 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$16947 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16948 VGND \$5637 \$411 \$5617 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$16949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16950 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16952 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16953 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16954 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16955 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16959 VPWR \$5638 VGND VPWR \$2908 VGND sky130_fd_sc_hd__clkbuf_1
X$16960 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16961 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16962 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16963 VPWR \$5653 VGND VPWR \$5638 VGND sky130_fd_sc_hd__clkbuf_1
X$16964 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16965 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16966 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16967 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16968 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16969 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16970 VPWR VGND sram_ro_addr[6] VPWR \$461 VGND sky130_fd_sc_hd__buf_2
X$16971 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16972 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16973 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16974 VGND \$470 \$481 \$387 \$491 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$16975 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16976 VPWR \$438 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$16977 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$16978 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16979 VPWR \$470 VGND VPWR \$438 VGND sky130_fd_sc_hd__clkbuf_1
X$16980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$16981 VPWR VGND \$428 VPWR \$439 \$374 \$462 VGND sky130_fd_sc_hd__a21oi_1
X$16982 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16983 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16984 VPWR \$462 VGND \$428 VPWR \$439 VGND sky130_fd_sc_hd__nor2_1
X$16985 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16986 VPWR \$439 \$382 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$16987 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$16988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16989 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16990 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16991 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16992 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$16993 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$16994 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$16995 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$16996 VGND \$455 \$428 \$471 \$492 \$482 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$16997 VPWR VGND VPWR \$471 \$440 VGND sky130_fd_sc_hd__inv_2
X$16998 VPWR \$472 VGND VPWR \$441 VGND sky130_fd_sc_hd__clkbuf_1
X$16999 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17000 VGND \$472 \$482 \$381 \$455 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$17001 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17002 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17003 VPWR \$483 VGND VPWR \$493 VGND sky130_fd_sc_hd__clkbuf_1
X$17004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17005 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17006 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17007 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17008 VPWR VGND \$443 \$293 \$182 \$505 \$429 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17011 VPWR VGND \$443 \$294 \$350 \$444 \$429 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17012 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17013 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17014 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17015 VGND \$463 \$239 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17016 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17017 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17018 VPWR VGND VPWR \$485 \$350 VGND sky130_fd_sc_hd__inv_2
X$17019 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17023 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17024 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17025 VPWR \$473 \$373 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17026 VPWR \$204 \$205 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17027 VPWR \$506 \$398 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17029 VGND \$463 \$241 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17030 VPWR \$456 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17031 VPWR \$465 VGND \$456 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$17032 VPWR VGND \$205 VPWR \$465 VGND sky130_fd_sc_hd__buf_2
X$17033 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17034 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17035 VGND \$206 \$430 \$241 \$445 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$17036 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17037 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17038 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17039 VGND \$206 \$486 \$196 \$494 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17040 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17041 VPWR VGND VPWR \$475 \$430 VGND sky130_fd_sc_hd__inv_2
X$17042 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17043 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17045 VPWR \$431 VGND \$320 \$464 VPWR VGND sky130_fd_sc_hd__or2_1
X$17046 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17048 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17049 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17050 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17051 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17055 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17056 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17057 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17058 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17061 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17062 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17063 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17064 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17066 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17067 VGND \$497 \$216 \$433 \$420 \$476 \$477 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$17068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17069 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17070 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17071 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17072 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17074 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17075 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17076 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17077 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17079 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17081 VPWR \$499 VGND VPWR \$221 \$326 \$489 \$347 VGND
+ sky130_fd_sc_hd__o22a_1
X$17082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17083 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17084 VPWR VGND VPWR \$489 \$399 VGND sky130_fd_sc_hd__inv_2
X$17085 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17087 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17088 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17089 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17090 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17092 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17093 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17094 VPWR VGND \$417 \$281 \$458 \$450 \$434 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17095 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17096 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17097 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17098 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17099 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17100 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17101 VGND \$206 \$478 \$466 \$467 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17102 VGND \$458 \$500 VPWR VPWR VGND sky130_fd_sc_hd__inv_8
X$17103 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17104 VGND \$467 \$289 \$478 \$479 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$17105 VGND \$206 \$459 \$246 \$501 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17106 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17107 VGND \$479 \$459 \$421 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17108 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17109 VGND \$206 \$436 \$246 \$460 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17112 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17113 VGND \$510 \$436 \$511 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17114 VGND \$206 \$480 \$246 \$468 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17115 VGND \$490 \$480 \$633 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17116 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17117 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17118 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17119 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17121 VPWR \$1606 \$451 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17122 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17123 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17124 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17125 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17126 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17127 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17128 VPWR \$457 \$394 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17129 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17131 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17133 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17134 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17135 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17136 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17137 VPWR VPWR VGND \$503 \$306 VGND sky130_fd_sc_hd__clkbuf_2
X$17138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17140 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17141 VPWR VGND \$301 \$386 \$211 \$469 \$306 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17142 VGND \$211 \$254 \$469 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$17143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17144 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17145 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17148 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17149 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17151 VPWR VGND sram_ro_addr[3] VPWR \$343 VGND sky130_fd_sc_hd__buf_2
X$17152 VGND \$371 \$387 \$401 \$308 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17153 VPWR VGND sram_ro_addr[4] VPWR \$350 VGND sky130_fd_sc_hd__buf_2
X$17154 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17155 VPWR VGND sram_ro_addr[5] VPWR \$373 VGND sky130_fd_sc_hd__buf_2
X$17156 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17158 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17160 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17161 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17162 VGND \$397 \$382 \$381 \$374 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$17163 VPWR \$359 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$17164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17166 VPWR \$375 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$17167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17168 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17169 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17170 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17171 VPWR \$376 VGND VPWR \$375 VGND sky130_fd_sc_hd__clkbuf_1
X$17172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17173 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17174 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17175 VPWR \$377 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$17176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17177 VPWR \$388 VGND VPWR \$377 VGND sky130_fd_sc_hd__clkbuf_1
X$17178 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17179 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17180 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17181 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17182 VGND \$655 \$194 \$237 \$331 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17183 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17186 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17187 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17190 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17191 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17192 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17193 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17194 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17195 VPWR VPWR VGND \$352 \$195 VGND sky130_fd_sc_hd__clkbuf_2
X$17196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17197 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17198 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17199 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17200 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17201 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17203 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17204 VPWR \$352 VGND \$325 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$17205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17206 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17207 VPWR \$273 VGND \$353 \$345 VPWR VGND sky130_fd_sc_hd__or2_1
X$17208 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17209 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17210 VPWR VGND \$204 \$354 \$346 \$361 \$205 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17211 VGND \$206 \$346 \$241 \$361 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$17212 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17213 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17214 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17217 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17218 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17219 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17220 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17221 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17222 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17223 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17224 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17225 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17226 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17228 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17231 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17232 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17233 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17234 VGND \$463 \$198 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17235 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17236 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17237 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17239 VGND \$365 \$355 \$356 \$188 \$420 \$295 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17240 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17241 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17242 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17243 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17244 VPWR \$366 VGND VPWR \$357 VGND sky130_fd_sc_hd__clkbuf_1
X$17245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17246 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17247 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17248 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17249 VPWR VGND \$384 \$424 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17250 VGND \$358 \$243 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17251 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17252 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17253 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17254 VGND \$206 \$348 \$243 \$367 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17255 VPWR VGND \$271 \$183 \$348 \$367 \$288 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17256 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17257 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17259 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17260 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17262 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17263 VGND \$278 \$363 \$456 \$379 \$385 \$391 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$17264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17265 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17266 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17267 VPWR VGND \$417 \$354 \$339 \$349 \$434 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17268 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17269 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17270 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17272 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17273 VPWR VGND \$339 \$385 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17277 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17279 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17280 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17282 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17284 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17285 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17287 VGND \$340 \$289 \$341 \$490 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$17288 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17291 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17292 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17293 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17294 VGND \$206 \$393 \$246 \$392 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17295 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17296 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17298 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17299 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17301 VPWR VGND \$291 \$386 \$394 \$395 \$292 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17302 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17303 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17304 VGND \$206 \$396 \$246 \$369 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17305 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17306 VPWR VPWR VGND \$369 VGND sky130_fd_sc_hd__conb_1
X$17307 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17308 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17309 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17310 VGND \$380 \$394 \$396 \$300 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17311 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17314 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17315 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17316 VPWR VGND serial_data_1 VPWR \$304 VGND sky130_fd_sc_hd__buf_2
X$17317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17318 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17320 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17322 VPWR VGND \$1704 VPWR debug_oeb VGND sky130_fd_sc_hd__clkbuf_4
X$17323 VPWR \$2424 VPWR VGND \$2537 \$2015 VGND sky130_fd_sc_hd__or2_2
X$17324 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17325 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17326 VPWR \$2657 VGND \$2608 \$2677 VPWR VGND sky130_fd_sc_hd__or2_1
X$17327 VPWR \$2656 \$2426 \$2676 VPWR VGND \$2657 \$2624 VGND
+ sky130_fd_sc_hd__or4_1
X$17328 VPWR \$2657 \$2435 VGND \$2697 VPWR \$2678 \$2712 VGND
+ sky130_fd_sc_hd__or4_2
X$17329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17330 VPWR \$2658 \$2513 \$2677 VPWR VGND \$2697 \$2638 VGND
+ sky130_fd_sc_hd__or4_1
X$17331 VPWR VGND VPWR \$2677 \$2698 VGND sky130_fd_sc_hd__inv_2
X$17332 VPWR \$2638 VGND \$2472 VPWR \$2659 VGND sky130_fd_sc_hd__nor2_1
X$17333 VPWR \$2697 VGND \$2511 VPWR \$2659 VGND sky130_fd_sc_hd__nor2_1
X$17334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17335 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17336 VPWR \$2521 VGND \$2659 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$17337 VPWR \$3431 \$2660 \$2712 VPWR VGND \$2512 \$2365 VGND
+ sky130_fd_sc_hd__or4_1
X$17338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17340 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17341 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17342 VPWR VPWR \$2741 VGND \$2514 \$2679 \$2699 VGND sky130_fd_sc_hd__o21ai_1
X$17343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17344 VPWR \$1963 VGND \$1960 \$2680 VPWR \$2661 VGND sky130_fd_sc_hd__o21ai_2
X$17345 VGND \$2699 \$2661 \$2758 \$2713 \$2514 \$2700 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$17346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17347 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17348 VPWR \$2715 VGND \$2354 \$2714 VPWR VGND sky130_fd_sc_hd__or2_1
X$17349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17350 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17351 VPWR VPWR \$2700 VGND \$2453 \$2716 \$2701 VGND sky130_fd_sc_hd__o21ai_1
X$17352 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17354 VPWR VGND \$2412 VPWR \$2640 \$2681 \$2716 VGND sky130_fd_sc_hd__a21oi_1
X$17355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17357 VPWR \$2662 VGND \$2488 \$2742 VPWR VGND sky130_fd_sc_hd__or2_1
X$17358 VPWR VGND VPWR \$2641 \$2662 VGND sky130_fd_sc_hd__inv_2
X$17359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17360 VPWR \$2717 VPWR VGND \$2681 \$2662 VGND sky130_fd_sc_hd__nand2_1
X$17361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17363 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17364 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17365 VGND \$2663 \$2683 \$2682 \$2441 \$2660 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$17366 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17367 VPWR \$2683 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17370 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17371 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17372 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17374 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17375 VPWR \$2323 \$2702 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17380 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17382 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17383 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17386 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17387 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17388 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17389 VPWR VGND VPWR \$2684 \$2558 VGND sky130_fd_sc_hd__inv_2
X$17390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17391 VPWR VGND \$2703 \$293 \$2704 \$2718 \$2705 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17392 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17394 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17397 VPWR \$2626 VGND VPWR \$2684 \$2355 \$2644 \$923 VGND
+ sky130_fd_sc_hd__o22a_1
X$17398 VPWR \$2297 \$2704 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17399 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17401 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17402 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17403 VGND \$2706 \$2735 \$1256 \$2525 \$2458 \$2597 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17404 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17405 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17406 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17407 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17408 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17409 VPWR \$2720 VGND VPWR \$1007 \$2724 \$2719 \$2316 VGND
+ sky130_fd_sc_hd__o22a_1
X$17410 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17412 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17413 VPWR VGND VPWR \$2687 \$2721 \$2706 \$2723 \$2722 VGND
+ sky130_fd_sc_hd__and4_1
X$17414 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17415 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17416 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17417 VPWR \$2598 VGND VPWR \$2664 \$2665 \$2123 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$17418 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17419 VPWR \$2685 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17420 VPWR \$2560 VGND VPWR \$2685 \$2665 \$2297 \$2688 VGND
+ sky130_fd_sc_hd__o22a_1
X$17421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17422 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17424 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17426 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17427 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17428 VPWR \$2686 VGND VPWR \$687 \$2045 \$1240 \$1955 VGND
+ sky130_fd_sc_hd__o22a_1
X$17429 VPWR \$1283 VGND VPWR \$2667 \$1571 VGND sky130_fd_sc_hd__or2_4
X$17430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17431 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17432 VPWR VPWR VGND \$2725 \$2346 VGND sky130_fd_sc_hd__clkbuf_2
X$17433 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17436 VGND \$2707 \$2645 \$2327 \$2113 \$1845 \$2666 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17438 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17439 VPWR VGND VPWR \$2584 \$2727 \$2689 \$2707 \$2726 VGND
+ sky130_fd_sc_hd__and4_1
X$17440 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17443 VGND \$2374 \$2647 \$2667 \$927 \$2668 \$2648 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$17444 VPWR VGND VPWR \$387 \$2668 VGND sky130_fd_sc_hd__inv_4
X$17445 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17447 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17448 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17449 VGND \$2689 \$2626 \$1481 \$1198 \$2386 \$2708 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17450 VPWR \$2690 VGND VPWR \$2286 \$1966 \$2518 \$1951 VGND
+ sky130_fd_sc_hd__o22a_1
X$17451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17452 VGND \$2828 \$2690 \$2708 \$2043 \$1914 \$2603 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17453 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17454 VPWR \$2604 VGND VPWR \$2669 \$2670 \$1481 \$2646 VGND
+ sky130_fd_sc_hd__o22a_1
X$17455 VGND \$2568 \$2728 \$2691 \$2544 \$2545 \$2708 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17456 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17457 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17458 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17459 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17460 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17463 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17464 VGND \$2692 \$2650 \$2033 \$2065 \$2046 \$2671 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$17465 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17466 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17468 VGND \$2617 \$2927 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$17469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17470 VPWR \$2693 VPWR VGND \$1449 \$1360 \$1705 VGND sky130_fd_sc_hd__or3_1
X$17471 VGND \$2693 \$2830 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$17472 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17473 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17475 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17477 VGND \$2618 \$2651 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$17478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17479 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17480 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17481 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17482 VPWR \$2652 VGND \$2386 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$17483 VPWR VGND VPWR \$2708 \$2709 VGND sky130_fd_sc_hd__inv_2
X$17484 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17485 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17486 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17487 VPWR VGND \$2634 VPWR \$2652 VGND sky130_fd_sc_hd__clkbuf_4
X$17488 VPWR VGND \$2633 \$1594 \$2709 \$2736 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17489 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17491 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17492 VPWR VGND \$2633 \$1179 \$2635 \$2636 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17493 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17494 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17495 VPWR VGND VPWR \$2633 \$2634 VGND sky130_fd_sc_hd__inv_2
X$17496 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17497 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17498 VGND \$1152 \$2653 \$2450 \$2695 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17500 VPWR VGND \$2694 \$386 \$2653 \$2695 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17502 VPWR VGND \$2694 \$1594 \$2637 \$2654 \$2672 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17504 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17506 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17507 VPWR VGND \$2729 \$1803 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17509 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17510 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17511 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17512 VPWR \$2503 \$2710 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17513 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17514 VPWR VGND \$2730 \$1594 \$2710 \$2655 \$2711 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17516 VGND \$1874 \$2232 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17518 VGND \$1152 \$2696 \$2232 \$2673 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17519 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17520 VPWR \$2671 \$2696 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$17521 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17524 VPWR VGND spimemio_flash_io0_di VPWR \$310 VGND sky130_fd_sc_hd__buf_2
X$17525 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17526 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17527 VPWR \$1395 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17528 VPWR \$1395 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17529 VPWR spimemio_flash_io0_do VPWR VGND \$1395 VGND sky130_fd_sc_hd__buf_4
X$17530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17531 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17532 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17533 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17534 VGND \$5519 \$4864 \$4733 \$2571 \$5536 \$4833 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_1
X$17535 VPWR VGND \$2571 VPWR \$4733 \$5517 \$5536 VGND sky130_fd_sc_hd__a21oi_1
X$17536 VPWR \$5536 VGND \$2571 VPWR \$4733 VGND sky130_fd_sc_hd__nor2_1
X$17537 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17540 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17541 VPWR VGND VPWR \$5470 \$5520 VGND sky130_fd_sc_hd__inv_2
X$17542 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17543 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17544 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17545 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17546 VPWR \$5529 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$17547 VPWR \$5530 VGND VPWR \$5529 VGND sky130_fd_sc_hd__clkbuf_1
X$17548 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17549 VPWR VGND \$5504 \$5537 \$5496 \$5522 \$1078 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17550 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17551 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17552 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17555 VPWR \$5544 VGND VPWR \$864 VGND sky130_fd_sc_hd__clkbuf_1
X$17556 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17557 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17559 VGND \$5270 \$5538 \$5532 \$5339 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$17560 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17561 VGND \$5538 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$17562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17563 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17564 VPWR VGND \$5192 \$354 \$5539 \$5552 \$4803 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17565 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17566 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17567 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17568 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17569 VPWR VGND \$5539 \$3674 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17572 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17573 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17574 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17576 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17577 VPWR VGND \$5229 \$184 \$5505 \$5524 \$5207 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17578 VGND \$2777 \$5546 \$4994 \$5534 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$17579 VGND \$2777 \$5526 \$4994 \$5535 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17580 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17581 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17582 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17583 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17584 VPWR VGND \$5540 \$3587 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17586 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17587 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17588 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17589 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17590 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17591 VPWR VGND VPWR \$4124 \$5541 VGND sky130_fd_sc_hd__inv_2
X$17592 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17593 VGND \$4761 \$5548 \$5369 \$5547 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17594 VPWR \$4600 \$5548 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17595 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17596 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17597 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17598 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17599 VGND \$4761 \$5500 \$5334 \$5514 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$17600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17601 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17603 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17604 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17605 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17606 VPWR VGND \$5345 \$1171 \$5501 \$5518 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17608 VGND \$4764 \$5528 \$5298 \$5549 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$17609 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17610 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17611 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17612 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17613 VGND \$5550 \$3711 \$5542 \$3924 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17614 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17615 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17617 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17619 VGND spimemio_flash_io0_oeb \$226 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$17620 VPWR \$5564 VGND VPWR \$5075 \$5439 \$1523 \$5448 VGND
+ sky130_fd_sc_hd__o22a_1
X$17621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17622 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17624 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17625 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17627 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17628 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17629 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17631 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17633 VGND \$5530 \$5537 \$4106 \$5555 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17634 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17635 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17636 VGND \$5565 \$5485 \$4106 \$5556 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17637 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17638 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17639 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17640 VPWR \$5545 VGND VPWR \$5557 VGND sky130_fd_sc_hd__clkbuf_1
X$17641 VGND \$5557 \$5531 \$5566 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17642 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17643 VGND \$5032 \$5558 \$5567 \$5533 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17644 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17645 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17646 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17647 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17648 VGND \$2777 \$5539 \$5165 \$5552 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17649 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17650 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17651 VPWR VGND \$5559 \$4774 \$5570 \$5569 \$5553 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17652 VPWR VPWR VGND \$4678 \$5553 VGND sky130_fd_sc_hd__clkbuf_2
X$17653 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17654 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17655 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17656 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17657 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17658 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17659 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17660 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17661 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17662 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17663 VPWR VGND \$5525 \$1171 \$5546 \$5534 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17664 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17665 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17666 VGND \$2777 \$5540 \$5367 \$5560 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17668 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17669 VPWR \$4559 \$5561 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17670 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17671 VPWR VGND \$5562 \$4774 \$5561 \$5571 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17672 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17674 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17675 VGND \$3952 \$5369 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17676 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17677 VPWR VGND \$5562 \$354 \$5548 \$5547 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17678 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17681 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17682 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17683 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17684 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17685 VGND \$3952 \$5334 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17686 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17687 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17688 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17689 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17690 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17691 VGND \$4764 \$5542 \$5298 \$5563 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17692 VGND \$4764 \$5572 \$5298 \$5554 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17693 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17694 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17695 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17696 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17697 VPWR VGND spimemio_flash_io2_di VPWR \$5726 VGND sky130_fd_sc_hd__buf_2
X$17698 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17699 VPWR \$5726 VGND VPWR \$5595 VGND sky130_fd_sc_hd__clkbuf_1
X$17700 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17701 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17702 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17703 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17705 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17707 VPWR \$5682 VGND \$5727 \$5147 VPWR VGND sky130_fd_sc_hd__or2_1
X$17708 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17709 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17710 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17711 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17712 VPWR VGND VPWR \$5699 \$5659 VGND sky130_fd_sc_hd__inv_2
X$17713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17714 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17715 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17716 VPWR \$5716 VGND VPWR \$5728 VGND sky130_fd_sc_hd__clkbuf_1
X$17717 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17719 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17721 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17722 VGND \$5708 \$5649 \$5729 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17723 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17724 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17725 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17726 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17727 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17729 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17730 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17731 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17732 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17733 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17734 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17735 VPWR VGND \$5559 \$3694 \$5718 \$5734 \$5553 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17736 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17737 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17738 VGND \$2777 \$5725 \$5165 \$5735 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17739 VPWR VGND \$5388 \$3711 \$5725 \$5735 \$5390 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17740 VPWR VGND VPWR \$5388 \$5390 VGND sky130_fd_sc_hd__inv_2
X$17741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17742 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17743 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17744 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17745 VGND \$2777 \$5720 \$5408 \$5719 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$17746 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17747 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17748 VGND \$2777 \$5711 \$4994 \$5736 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17749 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17750 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17751 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17752 VPWR VGND \$5498 \$3711 \$5703 \$5721 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17753 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17754 VGND \$4761 \$5712 \$5367 \$5737 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$17755 VPWR VGND \$5562 \$3711 \$5704 \$5713 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17756 VPWR VGND VPWR \$5498 \$5463 VGND sky130_fd_sc_hd__inv_2
X$17757 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17758 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17759 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17764 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17765 VPWR VGND \$5627 \$1171 \$5730 \$5738 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17766 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17767 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17769 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17770 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17773 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17774 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17775 VGND \$4764 \$5722 \$5334 \$5723 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17777 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17778 VPWR \$5739 VGND VPWR \$5707 \$4724 \$5731 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$17779 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17781 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17782 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17783 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17784 VPWR \$5740 VGND VPWR \$5695 \$4724 \$5732 \$5373 VGND
+ sky130_fd_sc_hd__o22a_1
X$17785 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17786 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17787 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17788 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17790 VPWR VGND \$5733 VPWR spimemio_flash_io2_do VGND
+ sky130_fd_sc_hd__clkbuf_4
X$17791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17792 VGND \$5302 \$5002 \$5755 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$17793 VPWR \$5439 \$5448 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$17794 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17795 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17796 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17797 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17798 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17799 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17800 VPWR \$5727 VPWR VGND \$5745 \$5468 \$5715 VGND sky130_fd_sc_hd__or3_1
X$17801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17802 VPWR \$5583 \$5679 VPWR \$5679 VGND \$5727 \$5727 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$17803 VGND \$5573 \$5699 \$5458 \$5727 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17804 VPWR VGND VPWR \$5679 \$5684 VGND sky130_fd_sc_hd__inv_2
X$17805 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17806 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17807 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17808 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17809 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17810 VPWR \$5761 VGND VPWR \$5746 VGND sky130_fd_sc_hd__clkbuf_1
X$17811 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17812 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17813 VGND \$5728 \$5610 \$5762 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17815 VPWR \$5763 VGND VPWR \$5747 VGND sky130_fd_sc_hd__clkbuf_1
X$17816 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17817 VGND \$5747 \$5748 \$5764 \$5551 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17818 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17819 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17820 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17825 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17826 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17827 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17828 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17829 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17831 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17832 VPWR VGND VPWR \$5559 \$5553 VGND sky130_fd_sc_hd__inv_2
X$17833 VGND \$2777 \$5718 \$5165 \$5734 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17834 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17835 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17836 VPWR VGND \$5750 \$3514 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17837 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17838 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17839 VPWR VGND VPWR \$5751 \$1755 VGND sky130_fd_sc_hd__inv_4
X$17840 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17842 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17843 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17845 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17846 VPWR VGND \$5525 \$184 \$5711 \$5736 \$5512 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17847 VPWR VGND VPWR \$5525 \$5512 VGND sky130_fd_sc_hd__inv_2
X$17848 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17850 VGND \$2777 \$5752 \$5367 \$5757 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17851 VPWR VGND \$5752 \$4107 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$17852 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17853 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17854 VPWR VGND \$5562 \$1171 \$5712 \$5737 \$5527 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17855 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17856 VPWR VGND \$5498 \$3694 \$5741 \$5766 \$5463 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17857 VGND \$4761 \$5741 \$5367 \$5766 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17858 VPWR \$1821 \$5741 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$17859 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17860 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17861 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17862 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17863 VGND \$5697 \$1925 mgmt_gpio_out[26] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$17864 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17865 VPWR VGND \$5627 \$3694 \$5758 \$5767 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17866 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17867 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17868 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17870 VPWR VGND \$5627 \$184 \$5759 \$5742 \$5589 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17872 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17873 VGND \$5698 \$1949 mgmt_gpio_out[30] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$17874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17875 VPWR VGND \$5345 \$3711 \$5760 \$5768 \$5323 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17876 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17877 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17878 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17879 VPWR \$5769 VGND VPWR \$4562 VGND sky130_fd_sc_hd__clkbuf_1
X$17880 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17881 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17882 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17883 VGND \$4764 \$5732 \$5298 \$5740 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17884 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17885 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17886 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17887 VPWR VGND VPWR \$5753 \$3063 VGND sky130_fd_sc_hd__inv_4
X$17888 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17889 VPWR VGND wb_dat_o[22] VPWR \$5024 VGND sky130_fd_sc_hd__buf_2
X$17890 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17891 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17892 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17893 VPWR \$5012 VGND VPWR \$4622 \$4508 \$1975 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$17894 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17895 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17896 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17897 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17898 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17899 VPWR \$5013 VPWR VGND \$5025 \$4942 \$4986 VGND sky130_fd_sc_hd__or3_1
X$17900 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17901 VGND \$5026 \$1979 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17902 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17903 VPWR \$4511 VPWR VGND \$1962 \$5027 VGND sky130_fd_sc_hd__or2_2
X$17904 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17905 VGND \$4006 \$4986 \$4917 \$4930 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$17906 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17907 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17908 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17909 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17910 VPWR \$5028 VGND \$4006 \$4623 VPWR VGND sky130_fd_sc_hd__or2_1
X$17911 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17912 VPWR VGND VPWR \$4800 \$5028 VGND sky130_fd_sc_hd__inv_2
X$17913 VPWR \$5015 VPWR VGND \$5028 \$5014 VGND sky130_fd_sc_hd__nand2_1
X$17914 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17915 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17916 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17917 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17918 VPWR VGND \$1979 VPWR \$4758 \$4953 VGND sky130_fd_sc_hd__nor2_2
X$17919 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17920 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17921 VPWR \$5017 \$5030 VPWR \$5029 VGND VGND sky130_fd_sc_hd__and2_1
X$17922 VPWR \$4779 VPWR VGND \$5031 \$5030 VGND sky130_fd_sc_hd__nand2_1
X$17923 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17924 VGND \$5018 \$1725 \$4933 \$5032 \$1452 \$5033 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$17925 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17926 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17928 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17929 VGND \$4374 \$4811 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$17930 VGND \$4761 \$4955 \$4811 \$4992 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17931 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17932 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17933 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17934 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17935 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17937 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17938 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17939 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17940 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17941 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17943 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17944 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17945 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17946 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17947 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17948 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17949 VGND \$4353 \$5020 \$4850 \$5019 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17950 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17951 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17952 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17953 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17954 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17955 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17957 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17958 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17959 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17960 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17961 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17962 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17963 VPWR VGND \$5044 \$354 \$5036 \$5041 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$17964 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17965 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17966 VPWR \$5021 VPWR \$5007 \$5134 \$3924 VGND \$3869 VGND
+ sky130_fd_sc_hd__a22oi_1
X$17967 VPWR VGND VPWR \$3629 \$5036 VGND sky130_fd_sc_hd__inv_2
X$17968 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17969 VGND \$4764 \$5009 \$5006 \$5037 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17970 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17971 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17972 VGND \$4764 \$4984 \$4828 \$4999 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$17973 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17975 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$17976 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17977 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17978 VGND \$5011 \$411 \$5038 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$17979 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17980 VGND \$5039 \$2862 mgmt_gpio_out[12] VPWR VPWR VGND
+ sky130_fd_sc_hd__ebufn_8
X$17981 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17982 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17983 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17984 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$17985 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$17986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17987 VPWR \$4986 VPWR VGND \$4916 \$4941 VGND sky130_fd_sc_hd__or2_2
X$17988 VGND \$3342 \$4986 \$4917 \$5025 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$17989 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$17990 VPWR \$3892 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$17991 VPWR \$5003 VGND \$3892 \$4916 VPWR VGND sky130_fd_sc_hd__or2_1
X$17992 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$17993 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$17994 VPWR \$4977 VGND \$4394 \$4942 VPWR VGND sky130_fd_sc_hd__or2_1
X$17995 VPWR \$4891 \$5027 \$4853 VPWR VGND \$4864 \$4733 VGND
+ sky130_fd_sc_hd__or4_1
X$17996 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$17997 VPWR VGND VPWR \$5040 \$4986 VGND sky130_fd_sc_hd__inv_2
X$17998 VPWR \$5042 VGND \$5027 \$4603 VPWR VGND sky130_fd_sc_hd__or2_1
X$17999 VGND \$5042 \$4673 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_8
X$18000 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18001 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18002 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18003 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18004 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18005 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18006 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18007 VPWR \$4738 VGND \$4895 VPWR \$1897 VGND sky130_fd_sc_hd__nor2_1
X$18008 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18009 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18010 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18011 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18012 VPWR \$5050 VGND \$4913 VPWR \$5031 VGND sky130_fd_sc_hd__or2b_1
X$18013 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18014 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18015 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18016 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18017 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18018 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18019 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18020 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18021 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18022 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18023 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18024 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18025 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18027 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18028 VPWR VGND VPWR \$2763 \$5071 VGND sky130_fd_sc_hd__inv_2
X$18029 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18030 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18031 VPWR VGND \$5043 VPWR \$4619 VGND sky130_fd_sc_hd__clkbuf_4
X$18032 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18033 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18034 VPWR \$4118 \$5053 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18035 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18036 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18037 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18038 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18039 VPWR VGND \$5044 \$3711 \$4981 \$4995 \$5035 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18040 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18041 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18042 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18043 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18045 VGND \$4764 \$5054 \$4850 \$5045 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18046 VPWR VGND VPWR \$3188 \$5054 VGND sky130_fd_sc_hd__inv_2
X$18047 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18048 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18049 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18050 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18051 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18053 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18054 VGND \$4764 \$5036 \$5006 \$5041 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18055 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18056 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18057 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18058 VPWR VGND \$5046 \$184 \$5009 \$5037 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18059 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18060 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18061 VPWR VGND \$5046 \$1594 \$5010 \$5022 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18062 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18063 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18064 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18065 VPWR VGND VPWR \$5068 \$1599 VGND sky130_fd_sc_hd__inv_4
X$18066 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18067 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18068 VGND \$3952 \$4828 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$18069 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18070 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18071 VGND \$2989 \$5039 \$4828 \$5047 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18072 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18073 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18074 VPWR \$5057 VGND VPWR \$5048 VGND sky130_fd_sc_hd__clkbuf_1
X$18075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18076 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18077 VPWR VGND wb_dat_o[23] VPWR \$5059 VGND sky130_fd_sc_hd__buf_2
X$18078 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18079 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18081 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18082 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18084 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18085 VPWR \$5026 VPWR VGND \$4930 \$4942 \$4986 VGND sky130_fd_sc_hd__or3_1
X$18086 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18087 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18088 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18089 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18090 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18091 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18092 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18093 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18094 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18096 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18097 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18098 VPWR \$5069 VGND \$4738 VPWR \$5061 VGND sky130_fd_sc_hd__nor2_1
X$18099 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18100 VPWR \$4676 \$5062 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18101 VPWR VGND VPWR \$4727 \$5078 VGND sky130_fd_sc_hd__inv_2
X$18102 VPWR VGND VPWR \$4954 \$5094 VGND sky130_fd_sc_hd__inv_2
X$18103 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18104 VPWR \$5050 VPWR VGND \$5063 \$5060 VGND sky130_fd_sc_hd__nand2_1
X$18105 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18106 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18107 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18108 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18109 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18110 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18112 VPWR VGND \$4701 \$293 \$5051 \$5070 \$4677 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18113 VPWR VGND VPWR \$4701 \$4677 VGND sky130_fd_sc_hd__inv_2
X$18114 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18115 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18116 VPWR VGND \$5051 \$2522 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$18117 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18118 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18119 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18120 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18121 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18122 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18123 VPWR VGND VPWR \$3262 \$5064 VGND sky130_fd_sc_hd__inv_2
X$18124 VGND \$4761 \$5071 \$4813 \$5065 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18125 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18126 VPWR \$1466 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18127 VPWR \$5119 VGND \$1466 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$18128 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18129 VPWR VGND \$5086 \$1594 \$5052 \$5072 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18130 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18131 VPWR VGND VPWR \$3722 \$5052 VGND sky130_fd_sc_hd__inv_2
X$18132 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18133 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18134 VPWR VGND \$5086 \$4023 \$5053 \$5082 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18135 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18136 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18138 VPWR VGND VPWR \$3536 \$5066 VGND sky130_fd_sc_hd__inv_2
X$18139 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18140 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18141 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18142 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18145 VPWR \$3601 \$5067 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18146 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18147 VGND \$3952 \$4850 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$18148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18149 VPWR VGND \$5005 \$184 \$5054 \$5045 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18150 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18151 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18154 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18155 VGND \$4764 \$5073 \$4765 \$5055 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18156 VPWR VGND VPWR \$5073 \$3036 VGND sky130_fd_sc_hd__inv_4
X$18157 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18158 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18159 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18161 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18162 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18163 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18165 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18166 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18167 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18168 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18170 VGND \$5074 \$5068 \$4774 \$4686 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18172 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18173 VPWR VGND \$4650 \$411 \$5038 \$5056 \$4659 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18174 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18175 VGND \$2989 \$5038 \$4828 \$5056 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18177 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18178 VPWR \$2880 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18179 VPWR \$5048 VGND VPWR \$2880 VGND sky130_fd_sc_hd__clkbuf_1
X$18180 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18181 VPWR VGND mgmt_gpio_oeb[15] VPWR \$5057 VGND sky130_fd_sc_hd__buf_2
X$18182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18183 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18184 VPWR VGND wb_dat_o[24] VPWR \$5075 VGND sky130_fd_sc_hd__buf_2
X$18185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18186 VPWR \$5104 VGND VPWR \$4776 \$5076 \$1523 \$5077 VGND
+ sky130_fd_sc_hd__o22a_1
X$18187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18189 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18191 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18192 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18193 VGND \$5089 \$3440 \$4853 VPWR VPWR VGND sky130_fd_sc_hd__nor2_4
X$18194 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18195 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18196 VPWR \$5090 VGND \$1963 \$5148 VPWR VGND sky130_fd_sc_hd__or2_1
X$18197 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18198 VPWR \$5060 VGND \$5090 \$4476 VPWR VGND sky130_fd_sc_hd__or2_1
X$18199 VPWR \$3858 \$5111 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18200 VPWR \$5078 VPWR VGND \$4698 \$1998 \$4603 VGND sky130_fd_sc_hd__or3_1
X$18201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18202 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18203 VPWR \$4503 \$4777 \$4772 VGND VPWR \$5091 VGND sky130_fd_sc_hd__or3b_2
X$18204 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18205 VPWR \$5092 VGND \$4772 VPWR \$4569 VGND sky130_fd_sc_hd__nor2_1
X$18206 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18207 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18208 VPWR VGND \$4953 VPWR \$5093 VGND sky130_fd_sc_hd__buf_2
X$18209 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18210 VPWR VPWR \$1998 VGND \$4895 \$5061 \$5141 VGND sky130_fd_sc_hd__o21ai_1
X$18211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18212 VPWR \$5062 VGND \$2511 \$4953 VPWR VGND sky130_fd_sc_hd__or2_1
X$18213 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18214 VPWR \$5094 VGND \$2472 \$4953 VPWR VGND sky130_fd_sc_hd__or2_1
X$18215 VPWR \$5069 \$5095 VPWR \$5062 VGND VGND sky130_fd_sc_hd__and2_1
X$18216 VGND \$5078 \$5063 \$5094 \$5095 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$18217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18218 VPWR VPWR \$1897 VGND \$4953 \$4913 \$5079 VGND sky130_fd_sc_hd__o21ai_1
X$18219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18220 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18221 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18222 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18223 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18224 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18225 VGND \$2777 \$5051 \$4811 \$5070 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18226 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18227 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18228 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18229 VGND \$4761 \$5064 \$4811 \$5096 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18230 VPWR VPWR VGND \$4636 \$5080 VGND sky130_fd_sc_hd__clkbuf_2
X$18231 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18232 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18233 VPWR VGND \$5097 \$4023 \$5071 \$5065 \$5081 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18234 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18235 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18236 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18237 VGND \$4761 \$5052 \$4813 \$5072 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18238 VGND \$4761 \$5053 \$4813 \$5082 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18240 VPWR VGND \$5005 \$3711 \$5066 \$5128 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18241 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18242 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18243 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18244 VPWR VGND \$5005 \$542 \$5099 \$5098 \$4957 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18245 VPWR VGND VPWR \$5005 \$4957 VGND sky130_fd_sc_hd__inv_2
X$18246 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18247 VPWR \$4119 \$5083 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18249 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18250 VGND \$4353 \$5067 \$4850 \$5084 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18251 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18252 VPWR VGND \$4905 \$4023 \$5067 \$5084 \$5100 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18253 VPWR VGND VPWR \$3624 \$5085 VGND sky130_fd_sc_hd__inv_2
X$18254 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18255 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18256 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18257 VPWR VGND \$5108 \$2628 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$18258 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18259 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18260 VPWR VGND \$5086 \$542 \$5073 \$5055 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18261 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18262 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18264 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18265 VPWR \$3544 \$5087 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18268 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18269 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18270 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18272 VPWR VGND \$5046 \$354 \$5102 \$5101 \$4998 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18273 VPWR \$3828 \$5102 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18274 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18276 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18277 VPWR \$5103 VGND VPWR \$5074 VGND sky130_fd_sc_hd__clkbuf_1
X$18278 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18279 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18280 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18281 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18282 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18283 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18285 VPWR VGND VPWR \$4501 \$4492 VGND sky130_fd_sc_hd__inv_2
X$18286 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18287 VPWR \$5047 VGND VPWR \$5144 \$4492 \$5039 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$18288 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18291 VPWR VGND wb_dat_o[28] VPWR \$5280 VGND sky130_fd_sc_hd__buf_2
X$18292 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18293 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18294 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18295 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18296 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18297 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18299 VGND \$3892 \$4942 \$4930 \$5281 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$18300 VGND \$4394 \$5025 \$4916 \$5281 VPWR VPWR VGND sky130_fd_sc_hd__or3_4
X$18301 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18302 VPWR \$5245 VGND \$5274 VPWR \$4733 VGND sky130_fd_sc_hd__nor2_1
X$18303 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18304 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18305 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18306 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18307 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18308 VGND \$2571 \$3663 \$4673 VPWR VPWR VGND sky130_fd_sc_hd__nor2_4
X$18309 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18310 VPWR \$5290 VGND \$5106 \$5282 VPWR VGND sky130_fd_sc_hd__or2_1
X$18311 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18312 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18313 VPWR \$3663 \$5291 \$5290 VPWR VGND \$4777 \$5283 VGND
+ sky130_fd_sc_hd__or4_1
X$18314 VPWR \$5284 \$5258 VGND \$5269 VPWR \$5285 VGND sky130_fd_sc_hd__nor3_1
X$18315 VPWR \$5292 VPWR VGND \$5285 \$5202 \$5291 VGND sky130_fd_sc_hd__or3_1
X$18316 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18317 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18318 VPWR \$5284 \$5286 \$5293 VPWR VGND \$4520 \$5183 VGND
+ sky130_fd_sc_hd__or4_1
X$18319 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18320 VPWR \$5276 VGND \$5247 VPWR \$5294 VGND sky130_fd_sc_hd__nor2_1
X$18321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18322 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18323 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18324 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18325 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18326 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18328 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18329 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18330 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18331 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18332 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18334 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18335 VGND \$4761 \$5277 \$5165 \$5287 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18336 VGND \$4761 \$5250 \$4813 \$5295 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18337 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18338 VPWR VGND VPWR \$5086 \$5043 VGND sky130_fd_sc_hd__inv_2
X$18339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18343 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18344 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18345 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18347 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18350 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18351 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18354 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18355 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18357 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18358 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18364 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18365 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18366 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18367 VPWR \$3321 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18368 VGND \$5296 \$3321 \$5297 \$3438 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18371 VGND \$4764 \$5299 \$5298 \$5288 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18373 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18374 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18376 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18377 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18378 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18379 VPWR \$5289 VGND VPWR \$5278 VGND sky130_fd_sc_hd__clkbuf_1
X$18380 VPWR VGND mgmt_gpio_oeb[16] VPWR \$5289 VGND sky130_fd_sc_hd__buf_2
X$18381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18383 VPWR VGND wb_dat_o[29] VPWR \$5302 VGND sky130_fd_sc_hd__buf_2
X$18384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18385 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18386 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18387 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18388 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18389 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18391 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18392 VGND \$4942 \$5281 \$5282 \$4673 \$5025 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4b_1
X$18393 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18394 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18395 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18396 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18399 VGND \$5303 \$4268 \$4777 \$5304 \$3663 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$18400 VPWR \$5283 VPWR VGND \$4267 \$5284 \$5304 VGND sky130_fd_sc_hd__or3_1
X$18401 VGND \$5292 \$5275 \$3573 \$5303 VPWR VPWR VGND sky130_fd_sc_hd__nor3_4
X$18402 VGND \$5275 \$4311 \$5202 \$5285 \$5284 VPWR VPWR VGND
+ sky130_fd_sc_hd__or4_4
X$18403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18404 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18405 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18407 VPWR VGND VPWR \$5317 \$5176 VGND sky130_fd_sc_hd__inv_2
X$18408 VPWR \$5318 VGND \$5225 VPWR \$5317 VGND sky130_fd_sc_hd__nor2_1
X$18409 VPWR \$5301 \$5225 VPWR \$5305 VGND VGND sky130_fd_sc_hd__and2_1
X$18410 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18411 VPWR VGND VPWR \$5115 \$5301 VGND sky130_fd_sc_hd__inv_2
X$18412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18415 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18416 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18417 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18418 VPWR VGND VPWR \$5307 \$3364 VGND sky130_fd_sc_hd__inv_4
X$18419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18420 VPWR VGND VPWR \$5118 \$5080 VGND sky130_fd_sc_hd__inv_2
X$18421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18422 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18423 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18424 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18425 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18426 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18427 VPWR VGND \$5086 \$4774 \$5250 \$5295 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18428 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18429 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18430 VPWR VGND VPWR \$5364 \$4275 VGND sky130_fd_sc_hd__inv_4
X$18431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18432 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18433 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18434 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18436 VPWR \$4134 \$5308 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18439 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18440 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18441 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18442 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18443 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18444 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18445 VPWR VGND VPWR \$3404 \$5309 VGND sky130_fd_sc_hd__inv_2
X$18446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18447 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18448 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18449 VPWR VGND \$5086 \$354 \$5310 \$5320 \$5043 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18450 VPWR \$4029 \$5310 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18453 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18454 VPWR VGND \$5311 \$3527 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$18455 VPWR VGND \$5344 \$386 \$5311 \$5321 \$5312 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18456 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18457 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18458 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18459 VPWR VGND \$5312 VPWR \$4795 VGND sky130_fd_sc_hd__clkbuf_4
X$18460 VPWR VGND VPWR \$3518 \$5313 VGND sky130_fd_sc_hd__inv_2
X$18461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18463 VPWR VGND \$5323 VPWR \$4261 VGND sky130_fd_sc_hd__buf_2
X$18464 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18465 VGND \$4764 \$5297 \$5298 \$5314 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18466 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18467 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18468 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18469 VGND \$4764 \$5324 \$5298 \$5315 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18470 VGND \$4764 \$5325 \$4828 \$5356 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18471 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18472 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18473 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18474 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18475 VPWR VGND sram_ro_clk VPWR \$555 VGND sky130_fd_sc_hd__buf_2
X$18476 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18477 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18479 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18480 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18481 VPWR \$583 VGND VPWR \$351 VGND sky130_fd_sc_hd__clkbuf_1
X$18482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18483 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18484 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18485 VGND \$536 \$564 \$574 \$599 \$440 VPWR VPWR VGND
+ sky130_fd_sc_hd__a31o_1
X$18486 VPWR \$544 VGND VPWR \$565 VGND sky130_fd_sc_hd__clkbuf_1
X$18487 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18488 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18489 VPWR \$585 VGND \$440 VPWR \$492 VGND sky130_fd_sc_hd__nor2_1
X$18490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18491 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18492 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18493 VPWR \$586 VGND VPWR \$565 VGND sky130_fd_sc_hd__clkbuf_1
X$18494 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18495 VGND \$587 \$555 \$293 \$523 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18496 VGND \$463 \$237 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$18497 VPWR VGND VPWR \$556 \$555 VGND sky130_fd_sc_hd__inv_2
X$18498 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18500 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18501 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18502 VGND \$575 \$524 \$686 \$557 \$1103 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_4
X$18503 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18504 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18505 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18506 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18507 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18508 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18509 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18510 VGND \$516 \$547 \$196 \$559 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18511 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18512 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18513 VPWR \$523 VPWR VGND \$566 \$345 VGND sky130_fd_sc_hd__or2_2
X$18514 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18515 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18516 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18517 VGND \$589 \$527 \$420 \$566 \$556 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$18518 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18519 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18520 VPWR VGND \$567 \$183 \$528 \$548 \$568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18521 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18522 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18523 VPWR VGND \$567 \$281 \$569 \$549 \$568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18524 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18525 VPWR \$590 \$552 VPWR \$539 VGND \$1103 \$560 VGND
+ sky130_fd_sc_hd__o2bb2a_1
X$18526 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18527 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18528 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18529 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18531 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18532 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18533 VPWR VGND VPWR \$576 \$518 VGND sky130_fd_sc_hd__inv_2
X$18534 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18535 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18536 VPWR \$570 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18537 VGND \$577 \$348 \$570 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18538 VPWR VGND VPWR \$579 \$406 VGND sky130_fd_sc_hd__inv_2
X$18539 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18540 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18541 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18542 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18543 VPWR \$580 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18545 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18546 VGND \$581 \$560 \$300 \$188 \$262 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2a_2
X$18547 VGND \$206 \$550 \$435 \$561 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18548 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18549 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18550 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18551 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18552 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18553 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18554 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18555 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18556 VPWR VGND VPWR \$520 \$560 VGND sky130_fd_sc_hd__inv_4
X$18557 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18559 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18560 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18561 VGND \$206 \$591 \$541 \$582 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18564 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18566 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18567 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18568 VGND \$201 \$552 \$571 \$300 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18569 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18571 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18572 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18574 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18575 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18576 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18577 VGND \$629 \$597 \$387 \$596 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$18578 VGND \$481 \$598 \$597 \$439 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$18579 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18580 VPWR \$584 VPWR VGND \$564 \$598 VGND sky130_fd_sc_hd__nand2_1
X$18581 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18582 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18583 VGND \$408 \$598 \$564 \$235 \$599 \$584 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$18584 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18585 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18586 VGND \$613 \$492 \$381 \$600 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18587 VGND \$565 \$351 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$18588 VPWR \$614 VGND VPWR \$587 VGND sky130_fd_sc_hd__clkbuf_1
X$18589 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18590 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18591 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18592 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18593 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18594 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18595 VPWR \$545 \$525 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18596 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18597 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18598 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18599 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18600 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18601 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18602 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18603 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18604 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18605 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18606 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18607 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18608 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18609 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18610 VPWR VGND \$547 \$601 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$18611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18612 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18613 VPWR VGND \$602 \$200 \$603 \$625 \$674 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18614 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18615 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18616 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18617 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18618 VPWR VGND \$567 \$200 \$604 \$632 \$568 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18619 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18620 VPWR VGND VPWR \$567 \$568 VGND sky130_fd_sc_hd__inv_2
X$18621 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18622 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18623 VPWR \$616 \$569 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18624 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18625 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18626 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18627 VGND \$516 \$617 \$605 \$606 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18628 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18629 VPWR VGND \$627 \$200 \$608 \$618 \$607 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18631 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18633 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18634 VPWR \$609 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18635 VGND \$368 \$223 \$609 \$578 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18636 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18637 VPWR \$619 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18638 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18639 VGND \$305 \$296 \$580 \$531 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18640 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18641 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18642 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18643 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18644 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18645 VPWR VGND \$550 \$620 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$18646 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18647 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18649 VGND \$651 \$289 \$593 \$822 \$251 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$18650 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18652 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18653 VGND \$427 \$610 \$577 \$322 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18654 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18657 VGND \$551 \$289 \$562 \$594 \$611 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$18658 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18659 VGND \$582 \$289 \$591 \$595 \$612 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$18660 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18661 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18662 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18663 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18664 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18665 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18666 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18667 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18668 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18669 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18670 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18671 VPWR VGND wb_dat_o[12] VPWR \$4601 VGND sky130_fd_sc_hd__buf_2
X$18672 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18673 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18674 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18675 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18676 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18678 VPWR \$4548 VPWR VGND \$4474 \$2472 \$4510 VGND sky130_fd_sc_hd__or3_1
X$18679 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18680 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18681 VPWR \$4615 VPWR \$4419 VGND \$4305 \$4633 VGND sky130_fd_sc_hd__o21a_1
X$18682 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18683 VPWR \$4443 VGND \$4477 \$4602 VPWR VGND sky130_fd_sc_hd__or2_1
X$18684 VPWR \$4305 \$4576 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18685 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18686 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18687 VGND \$4596 \$4603 \$1962 \$4035 \$4616 \$4604 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_1
X$18688 VGND \$2214 \$4578 \$4512 \$4597 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$18689 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18690 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18691 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18692 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18693 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18694 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18695 VPWR \$4605 \$4617 VGND \$4665 VPWR \$4158 \$4269 VGND
+ sky130_fd_sc_hd__or4_2
X$18696 VGND \$4287 \$4581 \$4605 \$4665 VPWR VPWR \$4617 VGND
+ sky130_fd_sc_hd__or4b_1
X$18697 VPWR \$4519 VGND \$4580 \$4572 VPWR VGND sky130_fd_sc_hd__or2_1
X$18698 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18699 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18700 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18701 VPWR VGND \$4555 \$4023 \$4606 \$4618 \$4530 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18703 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18704 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18705 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18706 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18707 VGND \$4353 \$4598 \$3921 \$4607 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18708 VPWR VGND \$4270 \$3711 \$4598 \$4607 \$4272 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18709 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18710 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18711 VGND \$1406 \$795 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$18712 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18713 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18714 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18715 VPWR \$4619 VGND \$3019 \$1406 VPWR VGND sky130_fd_sc_hd__or2_1
X$18716 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18717 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18718 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18719 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18721 VPWR \$4608 VGND VPWR \$4559 \$2447 \$2522 \$3621 VGND
+ sky130_fd_sc_hd__o22a_1
X$18722 VGND \$3868 \$4608 \$4609 \$2474 \$3553 \$2685 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18723 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18724 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18725 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18726 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18727 VPWR \$4599 VGND VPWR \$4480 \$2614 \$3645 \$1561 VGND
+ sky130_fd_sc_hd__o22a_1
X$18728 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18729 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18730 VPWR VGND VPWR \$3866 \$4610 VGND sky130_fd_sc_hd__inv_2
X$18731 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18732 VPWR VGND \$4407 \$542 \$4591 \$4590 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18733 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18734 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18735 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18736 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18737 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18738 VGND \$4611 \$4294 \$1089 \$1625 \$3587 \$2632 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$18739 VGND \$4342 \$4612 \$2481 \$2330 \$2219 \$4625 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18740 VPWR \$4611 VGND \$2447 \$4600 VPWR VGND sky130_fd_sc_hd__or2_1
X$18741 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18742 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18743 VPWR \$1134 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$18744 VPWR \$4620 VGND VPWR \$4088 \$2229 \$1134 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$18745 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18746 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18747 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18749 VGND \$4353 \$4593 \$4427 \$4592 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18750 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18751 VGND \$2989 \$4594 \$4427 \$4595 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18752 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18753 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18754 VPWR \$4244 \$4613 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18755 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18756 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18757 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18758 VGND \$3869 \$2919 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$18759 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18760 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18761 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18762 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18764 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18765 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18766 VPWR VGND wb_dat_o[13] VPWR \$4622 VGND sky130_fd_sc_hd__buf_2
X$18767 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18768 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18769 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18770 VGND \$3854 \$4367 \$4632 \$4548 VPWR VPWR VGND sky130_fd_sc_hd__and3_1
X$18771 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18772 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18773 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18774 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18775 VPWR VGND VPWR \$4633 \$4602 VGND sky130_fd_sc_hd__inv_2
X$18776 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18777 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18779 VPWR \$4616 VPWR VGND \$3342 \$4035 \$4603 VGND sky130_fd_sc_hd__or3_1
X$18780 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18781 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18782 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18783 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18784 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18785 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18786 VGND \$2742 \$4517 \$4623 \$2996 \$4623 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22ai_2
X$18787 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18789 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18790 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18791 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18792 VPWR VGND \$4555 \$3711 \$4634 \$4647 \$4530 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18793 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18794 VGND \$2777 \$4606 \$4216 \$4618 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18795 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18796 VPWR \$3643 \$4606 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18797 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18798 VPWR \$4635 VGND \$3621 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$18799 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18800 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18801 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18802 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18803 VPWR \$4636 VGND \$3204 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$18804 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18805 VPWR \$4637 VGND \$3556 \$795 VPWR VGND sky130_fd_sc_hd__or2_1
X$18806 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18808 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18809 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18810 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18811 VPWR VGND VPWR \$2518 \$4624 VGND sky130_fd_sc_hd__inv_2
X$18812 VPWR \$4638 VGND \$2497 \$804 VPWR VGND sky130_fd_sc_hd__or2_1
X$18813 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18814 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18815 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18816 VPWR VGND VPWR \$3403 \$4648 VGND sky130_fd_sc_hd__inv_2
X$18817 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18818 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18819 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18820 VPWR VGND VPWR \$3794 \$4669 VGND sky130_fd_sc_hd__inv_2
X$18821 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18822 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18823 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18824 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18825 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18826 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18827 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18828 VGND \$3952 \$4424 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$18829 VGND \$3903 \$4639 \$4319 \$2162 \$1089 \$4278 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18830 VPWR \$4639 VGND VPWR \$3403 \$2497 \$4625 \$2667 VGND
+ sky130_fd_sc_hd__o22a_1
X$18831 VPWR \$4612 VGND VPWR \$4058 \$2229 \$4670 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$18832 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18833 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18834 VPWR \$4626 VGND VPWR \$4029 \$2229 \$3675 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$18835 VGND \$4356 \$4626 \$4600 \$2330 \$2219 \$4627 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18836 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18837 VGND \$4209 \$4620 \$4628 \$2330 \$2219 \$3677 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18838 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18839 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18840 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18841 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18842 VPWR \$4357 \$4358 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18843 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18845 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18846 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18847 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18848 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18850 VGND \$4492 \$345 \$4629 \$4239 \$2919 VPWR VPWR VGND
+ sky130_fd_sc_hd__a211o_4
X$18851 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18852 VGND \$2989 \$4564 \$4165 \$4640 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18853 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18854 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18855 VGND \$4621 \$542 \$4641 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18856 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18857 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18858 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18859 VPWR \$4630 VGND VPWR \$4631 VGND sky130_fd_sc_hd__clkbuf_1
X$18860 VPWR VGND mgmt_gpio_oeb[13] VPWR \$4630 VGND sky130_fd_sc_hd__buf_2
X$18861 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18862 VPWR VGND wb_dat_o[11] VPWR \$4538 VGND sky130_fd_sc_hd__buf_2
X$18863 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18864 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18865 VGND \$4393 \$3277 \$4539 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$18866 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18867 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18868 VGND \$4474 \$4567 \$4548 \$4441 VPWR \$3430 VPWR VGND
+ sky130_fd_sc_hd__o211ai_4
X$18869 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18870 VPWR \$2214 VGND \$4540 \$3975 VPWR \$4549 VGND sky130_fd_sc_hd__o21ai_2
X$18871 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18872 VPWR \$4540 VGND \$4511 VPWR \$4444 VGND sky130_fd_sc_hd__nor2_1
X$18873 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18874 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18875 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18876 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18877 VPWR \$4527 VGND \$4513 \$4577 VPWR VGND sky130_fd_sc_hd__or2_1
X$18878 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18879 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18880 VPWR \$4551 \$4446 \$4528 VPWR VGND \$4515 \$4550 VGND
+ sky130_fd_sc_hd__or4_1
X$18881 VPWR \$4569 VGND \$4478 \$4459 VPWR VGND sky130_fd_sc_hd__or2_1
X$18882 VPWR \$4551 VPWR VGND \$4267 \$4153 \$4326 VGND sky130_fd_sc_hd__or3_1
X$18883 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18884 VPWR \$4494 VPWR VGND \$4153 \$4570 \$4517 VGND sky130_fd_sc_hd__or3_1
X$18885 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18886 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18887 VPWR \$4518 VGND \$4521 \$4552 \$4571 VPWR \$4553 VGND
+ sky130_fd_sc_hd__nor4_1
X$18888 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18889 VGND \$4504 \$4541 \$4520 \$4552 VPWR VPWR \$4572 VGND
+ sky130_fd_sc_hd__or4b_1
X$18890 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18891 VPWR VGND VPWR \$4573 \$4541 VGND sky130_fd_sc_hd__inv_2
X$18892 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18893 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18894 VGND \$2777 \$4542 \$4216 \$4554 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18895 VPWR VGND \$4555 \$3694 \$4542 \$4554 \$4530 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18896 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18897 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18898 VGND \$4353 \$4531 \$3921 \$4532 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18899 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18900 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18901 VPWR VGND \$4270 \$4023 \$4543 \$4583 \$4272 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18902 VPWR \$3509 \$4598 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18903 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18904 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18905 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18906 VPWR VGND \$4405 \$1179 \$4534 \$4533 \$4376 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18907 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18908 VGND \$4353 \$4523 \$4406 \$4556 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$18909 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18910 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18911 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18912 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18913 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18914 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18915 VPWR \$4314 VGND VPWR \$4274 \$2986 \$4544 \$2667 VGND
+ sky130_fd_sc_hd__o22a_1
X$18916 VGND \$4341 \$4557 \$4315 \$2330 \$2219 \$4544 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18917 VGND \$2004 \$3129 \$3621 \$2667 \$4558 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_2
X$18918 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18919 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18920 VPWR VGND \$4407 \$1594 \$4546 \$4574 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18921 VPWR \$3446 \$4546 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18922 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18923 VGND \$4316 \$4545 \$4559 \$2330 \$2219 \$4560 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$18924 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18925 VGND \$4353 \$4535 \$4424 \$4536 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$18926 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18927 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18928 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18929 VPWR \$1521 \$4226 VPWR VGND VGND sky130_fd_sc_hd__inv_6
X$18930 VGND \$4561 \$1521 \$1676 \$2447 \$4562 \$3165 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$18931 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18932 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18933 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18934 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18935 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18936 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18937 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18938 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18939 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18940 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18941 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18942 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18943 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18944 VPWR VGND \$4303 \$354 \$4563 \$4587 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$18945 VPWR \$4279 \$4563 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$18946 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18947 VPWR VGND VPWR \$4303 \$4321 VGND sky130_fd_sc_hd__inv_2
X$18948 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18949 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18950 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18951 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18952 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18953 VGND \$4547 \$1171 \$4564 \$3869 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$18954 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18955 VPWR \$4502 VGND VPWR \$4621 \$4492 \$4167 \$4501 VGND
+ sky130_fd_sc_hd__o22a_1
X$18956 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18957 VPWR VGND VPWR \$4526 \$4565 VGND sky130_fd_sc_hd__inv_2
X$18958 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18959 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18960 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18961 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18962 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18963 VPWR \$4539 VGND VPWR \$4393 \$4508 \$1523 \$4509 VGND
+ sky130_fd_sc_hd__o22a_1
X$18964 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18965 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18966 VPWR \$4510 VPWR \$4567 VGND \$4211 \$2571 VGND sky130_fd_sc_hd__o21a_1
X$18967 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18968 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18969 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18970 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18971 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18972 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$18973 VGND \$4442 \$1963 \$4006 \$2552 \$4576 \$4476 VPWR VPWR VGND
+ sky130_fd_sc_hd__a311o_1
X$18974 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18975 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$18976 VPWR VGND \$4527 \$4568 \$4578 VPWR \$3664 \$4596 VGND
+ sky130_fd_sc_hd__or4b_2
X$18977 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18978 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18979 VPWR \$4603 \$4515 VGND \$4035 VPWR \$1979 VGND sky130_fd_sc_hd__nor3_1
X$18980 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18981 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18982 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18983 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18984 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$18985 VPWR \$4326 \$4579 \$4552 VPWR VGND \$4478 \$4570 VGND
+ sky130_fd_sc_hd__or4_1
X$18986 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18987 VPWR \$4553 \$4495 \$4517 VPWR VGND \$4579 \$4589 VGND
+ sky130_fd_sc_hd__or4_1
X$18988 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18989 VPWR \$4581 \$4413 VPWR \$4580 VGND \$4573 \$4582 VGND
+ sky130_fd_sc_hd__o211ai_1
X$18990 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$18991 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18992 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18993 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18994 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18995 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18996 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$18997 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$18998 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$18999 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19000 VPWR VGND VPWR \$4270 \$4272 VGND sky130_fd_sc_hd__inv_2
X$19001 VGND \$4353 \$4543 \$3921 \$4583 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19002 VPWR VGND VPWR \$2610 \$4543 VGND sky130_fd_sc_hd__inv_2
X$19003 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19004 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19005 VPWR VGND \$4405 \$3711 \$4523 \$4556 \$4376 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19006 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19007 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19008 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19009 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19010 VPWR \$4545 VGND VPWR \$3842 \$2229 \$1612 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$19011 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19012 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19013 VPWR \$4557 VGND VPWR \$4118 \$2229 \$1755 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$19014 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19015 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19016 VGND \$355 \$4584 \$1125 \$4585 \$1465 VPWR VPWR VGND
+ sky130_fd_sc_hd__o22a_4
X$19017 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19018 VGND \$4353 \$4546 \$4377 \$4574 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19019 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19020 VGND \$3845 \$4599 \$4560 \$2667 \$1676 \$3540 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19021 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19022 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19023 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19024 VGND \$4353 \$4591 \$4424 \$4590 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$19025 VGND \$1855 \$4591 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$19026 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19027 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19028 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19029 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19030 VPWR \$4561 VGND VPWR \$2846 \$2986 \$4481 \$2614 VGND
+ sky130_fd_sc_hd__o22a_1
X$19031 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19032 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19033 VGND \$4586 \$4562 \$2330 \$2219 \$4558 \$2903 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$19034 VPWR \$4586 VGND VPWR \$3036 \$2229 \$4584 \$844 VGND
+ sky130_fd_sc_hd__o22a_1
X$19035 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19036 VPWR VGND \$4357 \$411 \$4593 \$4592 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19037 VPWR VGND VPWR \$4086 \$4593 VGND sky130_fd_sc_hd__inv_2
X$19038 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19039 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19040 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19041 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19042 VPWR VGND \$4357 \$542 \$4594 \$4595 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19043 VPWR VGND VPWR \$2923 \$4594 VGND sky130_fd_sc_hd__inv_2
X$19044 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19045 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19046 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19047 VGND \$2989 \$4563 \$4165 \$4587 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19048 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19049 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19050 VPWR \$4588 VGND \$2117 \$2919 VPWR VGND sky130_fd_sc_hd__or2_1
X$19051 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19052 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19053 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19054 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19055 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19056 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19057 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19058 VPWR \$4565 VGND VPWR mgmt_gpio_in[13] VGND sky130_fd_sc_hd__clkbuf_1
X$19059 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19060 VPWR VGND debug_in VPWR \$2520 VGND sky130_fd_sc_hd__buf_2
X$19061 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19062 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19063 VPWR \$2570 VGND \$2424 \$1962 VPWR VGND sky130_fd_sc_hd__or2_1
X$19064 VPWR VGND VPWR \$2608 \$2570 VGND sky130_fd_sc_hd__inv_2
X$19065 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19066 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19067 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19068 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19069 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19070 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19071 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19072 VPWR \$2354 VGND \$2514 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$19073 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19074 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19075 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19076 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19077 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19078 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19079 VPWR \$2440 VGND \$2453 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$19080 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19081 VPWR \$2392 VGND \$2488 VPWR \$2552 VGND sky130_fd_sc_hd__nor2_1
X$19082 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19083 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19084 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19085 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19086 VPWR VGND \$1771 \$200 \$2555 \$2554 \$1815 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19087 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19088 VPWR \$2609 \$2555 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19089 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19090 VGND \$856 \$2557 \$2556 \$2572 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19091 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19092 VGND \$856 \$2558 \$1861 \$2573 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19093 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19094 VGND \$1816 \$2574 \$2593 \$2314 \$2355 \$2594 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19095 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19096 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19097 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19098 VGND \$2576 \$2595 \$2596 \$2031 \$1554 \$2485 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19099 VGND \$2578 \$2367 \$2576 \$2304 \$2734 \$2597 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_1
X$19100 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19101 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19102 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19103 VPWR \$2579 VGND VPWR \$702 \$2559 \$2611 \$2540 VGND
+ sky130_fd_sc_hd__o22a_1
X$19104 VGND \$2495 \$2579 \$2936 \$2750 \$2541 \$819 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19105 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19106 VGND \$2200 \$2598 \$2610 \$2544 \$2545 \$2088 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19107 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19108 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19109 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19111 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19112 VPWR \$2612 VGND VPWR \$2121 \$1729 \$1242 \$859 VGND
+ sky130_fd_sc_hd__o22a_1
X$19113 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19114 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19115 VPWR VGND VPWR \$2613 \$2580 \$1731 \$2563 \$2528 VGND
+ sky130_fd_sc_hd__and4_1
X$19116 VPWR \$1570 VGND VPWR \$2581 \$1420 VGND sky130_fd_sc_hd__or2_4
X$19117 VGND \$1734 \$575 \$2599 \$2497 \$1466 \$2600 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19118 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19119 VPWR VGND VPWR \$2583 \$1301 \$2769 \$2582 \$477 VGND
+ sky130_fd_sc_hd__and4_1
X$19120 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19121 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19122 VGND \$2585 \$2601 \$2602 \$2613 VPWR \$2221 VPWR VGND
+ sky130_fd_sc_hd__nand4_2
X$19123 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19124 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19125 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19127 VGND \$2589 \$2603 \$2005 \$2604 \$2504 VPWR VPWR VGND
+ sky130_fd_sc_hd__o211a_1
X$19128 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19129 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19130 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19131 VGND \$2606 \$321 \$2605 \$2386 \$859 \$1390 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19132 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19133 VPWR \$2569 VPWR VGND \$1438 \$1882 \$1679 VGND sky130_fd_sc_hd__or3_1
X$19134 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19135 VPWR \$1448 \$2617 \$1415 VPWR VGND \$1360 \$1705 VGND
+ sky130_fd_sc_hd__or4_1
X$19136 VGND \$2532 \$2616 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$19137 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19138 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19139 VPWR \$2618 VPWR VGND \$1449 \$1882 \$1705 VGND sky130_fd_sc_hd__or3_1
X$19140 VPWR \$2619 VPWR VGND \$1449 \$1360 \$1679 VGND sky130_fd_sc_hd__or3_1
X$19141 VGND \$2534 \$2545 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$19142 VPWR \$2605 \$2607 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19143 VGND \$1152 \$2607 \$2450 \$2592 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19144 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19145 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19146 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19147 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19148 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19149 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19150 VPWR \$2551 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19151 VPWR \$2620 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19152 VPWR \$2620 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19153 VPWR \$2620 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19154 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19156 VPWR \$2620 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19157 VPWR \$2620 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19158 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19159 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19160 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19161 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19162 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19163 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19164 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19165 VPWR debug_mode VPWR VGND \$1587 VGND sky130_fd_sc_hd__buf_4
X$19166 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19167 VPWR \$2622 \$2623 \$2608 VPWR VGND \$2435 \$2407 VGND
+ sky130_fd_sc_hd__or4_1
X$19168 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19169 VPWR \$2624 VGND \$2407 \$2638 VPWR VGND sky130_fd_sc_hd__or2_1
X$19170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19171 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19172 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19173 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19174 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19175 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19176 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19177 VGND \$2639 \$2224 \$2214 \$2640 \$2171 \$2412 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_1
X$19178 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19179 VPWR \$2642 VGND \$2440 \$2641 VPWR VGND sky130_fd_sc_hd__or2_1
X$19180 VPWR \$2643 VGND \$2641 \$2104 VPWR VGND sky130_fd_sc_hd__or2_1
X$19181 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19182 VPWR \$2553 VGND \$2488 VPWR \$2571 VGND sky130_fd_sc_hd__nor2_1
X$19183 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19184 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19185 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19186 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19187 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19188 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19189 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19190 VPWR \$2644 \$2490 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19191 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19192 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19193 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19194 VPWR \$2594 \$2557 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19195 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19196 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19197 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19199 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19200 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19201 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19202 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19203 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19204 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19205 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19206 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19207 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19208 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19209 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19210 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19211 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19212 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19213 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19214 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19215 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19216 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19217 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19218 VGND \$2602 \$2648 \$2625 \$1700 \$2581 \$2587 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111a_2
X$19219 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19220 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19221 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19222 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19224 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19225 VPWR \$2627 VGND VPWR \$1051 \$1114 \$2628 \$2375 VGND
+ sky130_fd_sc_hd__o22a_1
X$19226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19227 VPWR \$2629 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19228 VGND \$2631 \$2627 \$2629 \$1819 \$1198 \$2630 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19229 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19230 VPWR \$2632 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$19231 VGND \$2632 \$391 \$2649 \$2631 \$2606 VPWR VPWR VGND
+ sky130_fd_sc_hd__and4_2
X$19232 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19233 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19234 VPWR \$2650 VGND VPWR \$1320 \$1793 \$1225 \$1811 VGND
+ sky130_fd_sc_hd__o22a_1
X$19235 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19236 VGND \$2507 \$2665 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$19237 VGND \$2591 \$2688 VPWR VPWR VGND sky130_fd_sc_hd__buf_6
X$19238 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19239 VGND \$2619 \$2646 VPWR VPWR VGND sky130_fd_sc_hd__buf_8
X$19240 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19241 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19242 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19243 VPWR VGND \$2633 \$354 \$2607 \$2592 \$2634 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19244 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19246 VPWR VGND VPWR \$2400 \$2635 VGND sky130_fd_sc_hd__inv_2
X$19247 VGND \$1152 \$2635 \$2450 \$2636 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$19248 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19249 VPWR \$2603 \$2637 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19250 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19251 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19252 VGND \$1152 \$2637 \$2232 \$2654 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19253 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19254 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19255 VGND \$1152 \$2710 \$2232 \$2655 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19257 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19259 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19260 VPWR VGND wb_dat_o[8] VPWR \$4393 VGND sky130_fd_sc_hd__buf_2
X$19261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19262 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19263 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19264 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19265 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19266 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19267 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19268 VPWR VGND \$4074 VPWR \$3954 \$4395 \$4394 VGND sky130_fd_sc_hd__a21oi_1
X$19269 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19270 VPWR \$3954 VGND \$4113 \$4396 VPWR VGND sky130_fd_sc_hd__or2_1
X$19271 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19272 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19273 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19274 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19275 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19277 VPWR VGND VPWR \$4397 \$1963 VGND sky130_fd_sc_hd__inv_2
X$19278 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19280 VPWR \$4399 VGND \$4369 \$3808 VPWR VGND sky130_fd_sc_hd__or2_1
X$19281 VPWR \$4398 VPWR VGND \$4009 \$4371 VGND sky130_fd_sc_hd__nand2_1
X$19282 VPWR VGND VPWR \$4400 \$4371 VGND sky130_fd_sc_hd__inv_2
X$19283 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19284 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19285 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19286 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19287 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19288 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19289 VGND \$2777 \$4382 \$4216 \$4401 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19290 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19291 VGND \$4374 \$3813 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$19292 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19294 VPWR VGND \$4183 \$3694 \$4354 \$4360 \$4185 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19295 VPWR \$3564 \$4383 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19297 VGND \$4353 \$4403 \$3921 \$4402 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19299 VPWR VGND VPWR \$2515 \$4403 VGND sky130_fd_sc_hd__inv_2
X$19300 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19301 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19302 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19303 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19304 VPWR VGND \$4404 \$1817 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$19305 VPWR VGND \$4405 \$3732 \$4384 \$4385 \$4376 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19306 VGND \$4353 \$4384 \$4406 \$4385 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19307 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19308 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19309 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19310 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19311 VPWR VGND \$4407 \$4023 \$4386 \$4362 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19312 VPWR VGND VPWR \$1838 \$4386 VGND sky130_fd_sc_hd__inv_2
X$19313 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19314 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19315 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19316 VPWR \$4387 VGND VPWR \$3934 \$1810 \$3965 \$2375 VGND
+ sky130_fd_sc_hd__o22a_1
X$19317 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19318 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19319 VGND \$4387 \$3399 \$2162 \$1845 \$3967 \$2361 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$19320 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19321 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19322 VPWR VGND \$4407 \$184 \$4388 \$4416 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19323 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19324 VPWR VGND \$4407 \$411 \$4389 \$4378 \$4363 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19325 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19326 VPWR VGND VPWR \$2089 \$4390 VGND sky130_fd_sc_hd__inv_2
X$19327 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19329 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19330 VPWR VGND VPWR \$4258 \$4389 VGND sky130_fd_sc_hd__inv_2
X$19331 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19332 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19333 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19334 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19335 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19336 VGND \$4163 \$4408 \$1099 \$785 \$2220 \$1812 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19337 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19338 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19339 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19340 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19342 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19343 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19344 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19345 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19346 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19347 VPWR VGND VPWR \$2853 \$4409 VGND sky130_fd_sc_hd__inv_2
X$19348 VGND \$2989 \$4409 \$4165 \$4391 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19349 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19350 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19351 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19352 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19353 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19355 VPWR \$4380 VGND VPWR \$2862 VGND sky130_fd_sc_hd__clkbuf_1
X$19356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19357 VPWR VGND mgmt_gpio_oeb[12] VPWR \$4379 VGND sky130_fd_sc_hd__buf_2
X$19358 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19359 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19360 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19361 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19362 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19363 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19364 VPWR VPWR \$2742 VGND \$3742 \$4410 \$4430 VGND sky130_fd_sc_hd__o21ai_1
X$19365 VPWR \$4430 VGND \$4074 \$2741 VPWR VGND sky130_fd_sc_hd__or2_1
X$19366 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19367 VPWR \$4419 \$3680 \$4411 VPWR VGND \$4410 \$4395 VGND
+ sky130_fd_sc_hd__or4_1
X$19368 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19369 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19371 VPWR \$4195 VGND \$2224 VPWR \$4412 VGND sky130_fd_sc_hd__nor2_1
X$19372 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19373 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19374 VGND \$4432 \$2224 \$4512 \$4420 \$4400 \$4369 VPWR VPWR VGND
+ sky130_fd_sc_hd__a311o_1
X$19375 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19376 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19377 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19378 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19379 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19380 VGND \$2261 \$4421 \$4433 \$3507 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$19381 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19382 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19383 VGND \$3507 \$4413 \$4434 \$1922 VPWR VPWR VGND sky130_fd_sc_hd__mux2_4
X$19384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19385 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19386 VPWR VGND \$4234 \$3732 \$4382 \$4401 \$4224 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19387 VPWR VGND \$4234 \$4023 \$4383 \$4435 \$4224 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19388 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19389 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19390 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19391 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19393 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19394 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19395 VPWR VGND \$4270 \$1179 \$4403 \$4402 \$4272 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19396 VPWR \$3898 \$4414 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$19397 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19398 VGND \$4353 \$4404 \$3921 \$4415 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19399 VPWR VGND \$4405 \$3694 \$4404 \$4415 \$4376 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19400 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19401 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19402 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19403 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19404 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19405 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19406 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19407 VGND \$4302 \$4422 \$2763 \$785 \$2220 \$1838 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19408 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19409 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19410 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19411 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19412 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19413 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19415 VGND \$4423 \$3236 \$785 \$2220 \$3446 \$2902 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$19416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19417 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19418 VGND \$4353 \$4388 \$4424 \$4416 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19420 VPWR VGND \$4388 \$1812 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$19421 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19422 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$19423 VGND \$4417 \$4425 \$4123 \$785 \$2220 \$4258 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19424 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$19425 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19426 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19427 VPWR \$4426 VGND VPWR \$3188 \$1954 \$3478 \$2226 VGND
+ sky130_fd_sc_hd__o22a_1
X$19428 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19429 VGND \$4408 \$4426 \$4173 \$2358 \$2274 \$3480 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_1
X$19430 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19431 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19433 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19434 VPWR VGND \$4357 \$386 \$4390 \$4418 \$4358 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19435 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19436 VGND \$2989 \$4390 \$4427 \$4418 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$19437 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$19440 VPWR VGND \$4303 \$1594 \$4409 \$4391 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19441 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19442 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19443 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19444 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$19445 VPWR VGND \$4303 \$542 \$3319 \$4437 \$4321 VPWR VGND
+ sky130_fd_sc_hd__a22o_1
X$19446 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19447 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19448 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$19449 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19450 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$19451 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$19452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
.ENDS housekeeping

.SUBCKT sky130_fd_sc_hd__conb_1 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__buf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__o311a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o311a_2

.SUBCKT sky130_fd_sc_hd__a221o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a221o_2

.SUBCKT sky130_fd_sc_hd__o2bb2a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o2bb2a_2

.SUBCKT sky130_fd_sc_hd__nand4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nand4_2

.SUBCKT sky130_fd_sc_hd__o221a_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221a_4

.SUBCKT sky130_fd_sc_hd__nor2_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_8

.SUBCKT sky130_fd_sc_hd__or3b_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3b_4

.SUBCKT sky130_fd_sc_hd__dfstp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_2

.SUBCKT sky130_fd_sc_hd__a31oi_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a31oi_1

.SUBCKT sky130_fd_sc_hd__and2b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__and2b_1

.SUBCKT sky130_fd_sc_hd__dfstp_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_4

.SUBCKT sky130_fd_sc_hd__a22o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22o_2

.SUBCKT sky130_fd_sc_hd__dfrtn_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtn_1

.SUBCKT sky130_fd_sc_hd__and3b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__and3b_1

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkdlybuf4s25_1

.SUBCKT sky130_fd_sc_hd__nor3_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3_2

.SUBCKT sky130_fd_sc_hd__or4b_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4b_4

.SUBCKT sky130_fd_sc_hd__o21ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ai_4

.SUBCKT sky130_fd_sc_hd__o211ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211ai_2

.SUBCKT sky130_fd_sc_hd__a2111o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a2111o_1

.SUBCKT sky130_fd_sc_hd__a311oi_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a311oi_2

.SUBCKT sky130_fd_sc_hd__nand2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__o2111a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111a_2

.SUBCKT sky130_fd_sc_hd__a2111o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a2111o_2

.SUBCKT sky130_fd_sc_hd__o2111ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111ai_2

.SUBCKT sky130_fd_sc_hd__o31a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o31a_1

.SUBCKT sky130_fd_sc_hd__o211ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211ai_4

.SUBCKT sky130_fd_sc_hd__o2111ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111ai_1

.SUBCKT sky130_fd_sc_hd__o2111ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111ai_4

.SUBCKT sky130_fd_sc_hd__nor4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nor4_2

.SUBCKT sky130_fd_sc_hd__o221ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221ai_2

.SUBCKT sky130_fd_sc_hd__o221ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221ai_1

.SUBCKT sky130_fd_sc_hd__o311a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o311a_1

.SUBCKT sky130_fd_sc_hd__o22ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22ai_2

.SUBCKT sky130_fd_sc_hd__and4bb_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__and4bb_1

.SUBCKT sky130_fd_sc_hd__o22ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22ai_4

.SUBCKT sky130_fd_sc_hd__a41o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a41o_1

.SUBCKT sky130_fd_sc_hd__a311oi_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a311oi_1

.SUBCKT sky130_fd_sc_hd__nor4_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nor4_1

.SUBCKT sky130_fd_sc_hd__nor2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_2

.SUBCKT sky130_fd_sc_hd__or3b_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3b_2

.SUBCKT sky130_fd_sc_hd__o21ba_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ba_1

.SUBCKT sky130_fd_sc_hd__o21bai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21bai_1

.SUBCKT sky130_fd_sc_hd__a41o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a41o_2

.SUBCKT sky130_fd_sc_hd__a21o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21o_2

.SUBCKT sky130_fd_sc_hd__clkbuf_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_8

.SUBCKT sky130_fd_sc_hd__clkinvlp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinvlp_2

.SUBCKT sky130_fd_sc_hd__nor3_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3_1

.SUBCKT sky130_fd_sc_hd__a21bo_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21bo_2

.SUBCKT sky130_fd_sc_hd__a21bo_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21bo_1

.SUBCKT sky130_fd_sc_hd__nand4bb_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nand4bb_1

.SUBCKT sky130_fd_sc_hd__o32a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o32a_1

.SUBCKT sky130_fd_sc_hd__o21a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21a_1

.SUBCKT sky130_fd_sc_hd__o31ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o31ai_4

.SUBCKT sky130_fd_sc_hd__nand3b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nand3b_1

.SUBCKT sky130_fd_sc_hd__a32o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a32o_2

.SUBCKT sky130_fd_sc_hd__o21ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ai_2

.SUBCKT sky130_fd_sc_hd__buf_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_8

.SUBCKT sky130_fd_sc_hd__or4bb_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4bb_1

.SUBCKT sky130_fd_sc_hd__or4bb_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4bb_4

.SUBCKT sky130_fd_sc_hd__nand4_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nand4_1

.SUBCKT sky130_fd_sc_hd__or3_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3_4

.SUBCKT sky130_fd_sc_hd__or3b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3b_1

.SUBCKT sky130_fd_sc_hd__nor3_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3_4

.SUBCKT sky130_fd_sc_hd__nor2_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_4

.SUBCKT sky130_fd_sc_hd__nand2_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_4

.SUBCKT sky130_fd_sc_hd__or2b_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2b_2

.SUBCKT sky130_fd_sc_hd__a311o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a311o_1

.SUBCKT sky130_fd_sc_hd__and4b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__and4b_1

.SUBCKT sky130_fd_sc_hd__o211a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211a_2

.SUBCKT sky130_fd_sc_hd__a32o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a32o_1

.SUBCKT sky130_fd_sc_hd__or2b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2b_1

.SUBCKT sky130_fd_sc_hd__nand2_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_8

.SUBCKT sky130_fd_sc_hd__or4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4_2

.SUBCKT sky130_fd_sc_hd__o22ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22ai_1

.SUBCKT sky130_fd_sc_hd__or4_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4_1

.SUBCKT sky130_fd_sc_hd__a21oi_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21oi_1

.SUBCKT sky130_fd_sc_hd__inv_12 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_12

.SUBCKT sky130_fd_sc_hd__and2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__and2_1

.SUBCKT sky130_fd_sc_hd__a221o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a221o_1

.SUBCKT sky130_fd_sc_hd__mux2_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_8

.SUBCKT sky130_fd_sc_hd__or4b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4b_1

.SUBCKT sky130_fd_sc_hd__o211ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211ai_1

.SUBCKT sky130_fd_sc_hd__or4b_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4b_2

.SUBCKT sky130_fd_sc_hd__o221ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221ai_4

.SUBCKT sky130_fd_sc_hd__o21ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ai_1

.SUBCKT sky130_fd_sc_hd__or3_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3_1

.SUBCKT sky130_fd_sc_hd__o32a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o32a_2

.SUBCKT sky130_fd_sc_hd__dfxtp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__dfxtp_1

.SUBCKT sky130_fd_sc_hd__a31o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a31o_1

.SUBCKT sky130_fd_sc_hd__a211o_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a211o_4

.SUBCKT sky130_fd_sc_hd__or2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2_2

.SUBCKT sky130_fd_sc_hd__nand2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_1

.SUBCKT sky130_fd_sc_hd__nand4b_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nand4b_4

.SUBCKT sky130_fd_sc_hd__and3_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__and3_2

.SUBCKT sky130_fd_sc_hd__and3_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__and3_1

.SUBCKT sky130_fd_sc_hd__o2111a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111a_1

.SUBCKT sky130_fd_sc_hd__o22a_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22a_4

.SUBCKT sky130_fd_sc_hd__and3_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__and3_4

.SUBCKT sky130_fd_sc_hd__mux2_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_4

.SUBCKT sky130_fd_sc_hd__inv_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_8

.SUBCKT sky130_fd_sc_hd__clkinv_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_8

.SUBCKT sky130_fd_sc_hd__mux2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_2

.SUBCKT sky130_fd_sc_hd__ebufn_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__ebufn_2

.SUBCKT sky130_fd_sc_hd__a22oi_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22oi_1

.SUBCKT sky130_fd_sc_hd__inv_6 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_6

.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__dlymetal6s2s_1

.SUBCKT sky130_fd_sc_hd__a22oi_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22oi_4

.SUBCKT sky130_fd_sc_hd__inv_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_4

.SUBCKT sky130_fd_sc_hd__ebufn_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__ebufn_8

.SUBCKT sky130_fd_sc_hd__mux2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__o2bb2a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o2bb2a_1

.SUBCKT sky130_fd_sc_hd__dfrtp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_2

.SUBCKT sky130_fd_sc_hd__buf_12 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_12

.SUBCKT sky130_fd_sc_hd__nand3_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nand3_4

.SUBCKT sky130_fd_sc_hd__clkbuf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__nor2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_1

.SUBCKT sky130_fd_sc_hd__a2bb2o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a2bb2o_1

.SUBCKT sky130_fd_sc_hd__a21o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21o_1

.SUBCKT sky130_fd_sc_hd__clkinv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_2

.SUBCKT sky130_fd_sc_hd__and4_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__and4_1

.SUBCKT sky130_fd_sc_hd__clkbuf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__or3_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3_2

.SUBCKT sky130_fd_sc_hd__or4_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4_4

.SUBCKT sky130_fd_sc_hd__o211a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211a_1

.SUBCKT sky130_fd_sc_hd__clkbuf_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_4

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 nc_1 nc_2
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__decap_4 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__buf_6 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_6

.SUBCKT sky130_fd_sc_hd__buf_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_4

.SUBCKT sky130_fd_sc_hd__a211o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a211o_1

.SUBCKT sky130_fd_sc_hd__clkbuf_16 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_16

.SUBCKT sky130_fd_sc_hd__o221a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221a_2

.SUBCKT sky130_fd_sc_hd__nand4_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__nand4_4

.SUBCKT sky130_fd_sc_hd__o221a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221a_1

.SUBCKT sky130_fd_sc_hd__and4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__and4_2

.SUBCKT sky130_fd_sc_hd__fill_2 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__diode_2 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__or2_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2_4

.SUBCKT sky130_fd_sc_hd__dfrtp_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_4

.SUBCKT sky130_fd_sc_hd__decap_6 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__o22a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22a_1

.SUBCKT sky130_fd_sc_hd__clkinv_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_4

.SUBCKT sky130_fd_sc_hd__inv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__fill_1 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__o22a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22a_2

.SUBCKT sky130_fd_sc_hd__decap_8 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__dfrtp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_1

.SUBCKT sky130_fd_sc_hd__or2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2_1

.SUBCKT sky130_fd_sc_hd__decap_3 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__a22o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22o_1

.SUBCKT sky130_fd_sc_hd__dfstp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_1

.SUBCKT sky130_fd_sc_hd__buf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__decap_12 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_12
