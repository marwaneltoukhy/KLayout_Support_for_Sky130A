*
*  /home/marwan/ef/klayout_lvs/lvs/test_cases/mgmt_protect/mgmt_protect.spice : SPICE netlist translated from the VERILOG netlist : /home/marwan/ef/caravel/verilog/gl/mgmt_protect.v
*                                                                               on the 2021-12-22 17:56:37.361845
*
***************************************************************************************************************************************************************************************

.INCLUDE sky130_fd_sc_hd.spice 

.GLOBAL VDD VSS

.SUBCKT MGMT_PROTECT CARAVEL_CLK CARAVEL_CLK2 CARAVEL_RSTN MPRJ_ACK_I_CORE MPRJ_ACK_I_USER MPRJ_CYC_O_CORE MPRJ_CYC_O_USER MPRJ_IENA_WB MPRJ_STB_O_CORE MPRJ_STB_O_USER MPRJ_WE_O_CORE MPRJ_WE_O_USER USER1_VCC_POWERGOOD USER1_VDD_POWERGOOD USER2_VCC_POWERGOOD USER2_VDD_POWERGOOD USER_CLOCK USER_CLOCK2 USER_RESET VCCD VCCD1 VCCD2 VDDA1 VDDA2 VSSA1 VSSA2 VSSD VSSD1 VSSD2 LA_DATA_IN_CORE[0] LA_DATA_IN_CORE[1] LA_DATA_IN_CORE[2] LA_DATA_IN_CORE[3] LA_DATA_IN_CORE[4] LA_DATA_IN_CORE[5] LA_DATA_IN_CORE[6] LA_DATA_IN_CORE[7] LA_DATA_IN_CORE[8] LA_DATA_IN_CORE[9] LA_DATA_IN_CORE[10] LA_DATA_IN_CORE[11] LA_DATA_IN_CORE[12] LA_DATA_IN_CORE[13] LA_DATA_IN_CORE[14] LA_DATA_IN_CORE[15] LA_DATA_IN_CORE[16] LA_DATA_IN_CORE[17] LA_DATA_IN_CORE[18] LA_DATA_IN_CORE[19] LA_DATA_IN_CORE[20] LA_DATA_IN_CORE[21] LA_DATA_IN_CORE[22] LA_DATA_IN_CORE[23] LA_DATA_IN_CORE[24] LA_DATA_IN_CORE[25] LA_DATA_IN_CORE[26] LA_DATA_IN_CORE[27] LA_DATA_IN_CORE[28] LA_DATA_IN_CORE[29] LA_DATA_IN_CORE[30] LA_DATA_IN_CORE[31] LA_DATA_IN_CORE[32] LA_DATA_IN_CORE[33] LA_DATA_IN_CORE[34] LA_DATA_IN_CORE[35] LA_DATA_IN_CORE[36] LA_DATA_IN_CORE[37] LA_DATA_IN_CORE[38] LA_DATA_IN_CORE[39] LA_DATA_IN_CORE[40] LA_DATA_IN_CORE[41] LA_DATA_IN_CORE[42] LA_DATA_IN_CORE[43] LA_DATA_IN_CORE[44] LA_DATA_IN_CORE[45] LA_DATA_IN_CORE[46] LA_DATA_IN_CORE[47] LA_DATA_IN_CORE[48] LA_DATA_IN_CORE[49] LA_DATA_IN_CORE[50] LA_DATA_IN_CORE[51] LA_DATA_IN_CORE[52] LA_DATA_IN_CORE[53] LA_DATA_IN_CORE[54] LA_DATA_IN_CORE[55] LA_DATA_IN_CORE[56] LA_DATA_IN_CORE[57] LA_DATA_IN_CORE[58] LA_DATA_IN_CORE[59] LA_DATA_IN_CORE[60] LA_DATA_IN_CORE[61] LA_DATA_IN_CORE[62] LA_DATA_IN_CORE[63] LA_DATA_IN_CORE[64] LA_DATA_IN_CORE[65] LA_DATA_IN_CORE[66] LA_DATA_IN_CORE[67] LA_DATA_IN_CORE[68] LA_DATA_IN_CORE[69] LA_DATA_IN_CORE[70] LA_DATA_IN_CORE[71] LA_DATA_IN_CORE[72] LA_DATA_IN_CORE[73] LA_DATA_IN_CORE[74] LA_DATA_IN_CORE[75] LA_DATA_IN_CORE[76] LA_DATA_IN_CORE[77] LA_DATA_IN_CORE[78] LA_DATA_IN_CORE[79] LA_DATA_IN_CORE[80] LA_DATA_IN_CORE[81] LA_DATA_IN_CORE[82] LA_DATA_IN_CORE[83] LA_DATA_IN_CORE[84] LA_DATA_IN_CORE[85] LA_DATA_IN_CORE[86] LA_DATA_IN_CORE[87] LA_DATA_IN_CORE[88] LA_DATA_IN_CORE[89] LA_DATA_IN_CORE[90] LA_DATA_IN_CORE[91] LA_DATA_IN_CORE[92] LA_DATA_IN_CORE[93] LA_DATA_IN_CORE[94] LA_DATA_IN_CORE[95] LA_DATA_IN_CORE[96] LA_DATA_IN_CORE[97] LA_DATA_IN_CORE[98] LA_DATA_IN_CORE[99] LA_DATA_IN_CORE[100] LA_DATA_IN_CORE[101] LA_DATA_IN_CORE[102] LA_DATA_IN_CORE[103] LA_DATA_IN_CORE[104] LA_DATA_IN_CORE[105] LA_DATA_IN_CORE[106] LA_DATA_IN_CORE[107] LA_DATA_IN_CORE[108] LA_DATA_IN_CORE[109] LA_DATA_IN_CORE[110] LA_DATA_IN_CORE[111] LA_DATA_IN_CORE[112] LA_DATA_IN_CORE[113] LA_DATA_IN_CORE[114] LA_DATA_IN_CORE[115] LA_DATA_IN_CORE[116] LA_DATA_IN_CORE[117] LA_DATA_IN_CORE[118] LA_DATA_IN_CORE[119] LA_DATA_IN_CORE[120] LA_DATA_IN_CORE[121] LA_DATA_IN_CORE[122] LA_DATA_IN_CORE[123] LA_DATA_IN_CORE[124] LA_DATA_IN_CORE[125] LA_DATA_IN_CORE[126] LA_DATA_IN_CORE[127] LA_DATA_IN_MPRJ[0] LA_DATA_IN_MPRJ[1] LA_DATA_IN_MPRJ[2] LA_DATA_IN_MPRJ[3] LA_DATA_IN_MPRJ[4] LA_DATA_IN_MPRJ[5] LA_DATA_IN_MPRJ[6] LA_DATA_IN_MPRJ[7] LA_DATA_IN_MPRJ[8] LA_DATA_IN_MPRJ[9] LA_DATA_IN_MPRJ[10] LA_DATA_IN_MPRJ[11] LA_DATA_IN_MPRJ[12] LA_DATA_IN_MPRJ[13] LA_DATA_IN_MPRJ[14] LA_DATA_IN_MPRJ[15] LA_DATA_IN_MPRJ[16] LA_DATA_IN_MPRJ[17] LA_DATA_IN_MPRJ[18] LA_DATA_IN_MPRJ[19] LA_DATA_IN_MPRJ[20] LA_DATA_IN_MPRJ[21] LA_DATA_IN_MPRJ[22] LA_DATA_IN_MPRJ[23] LA_DATA_IN_MPRJ[24] LA_DATA_IN_MPRJ[25] LA_DATA_IN_MPRJ[26] LA_DATA_IN_MPRJ[27] LA_DATA_IN_MPRJ[28] LA_DATA_IN_MPRJ[29] LA_DATA_IN_MPRJ[30] LA_DATA_IN_MPRJ[31] LA_DATA_IN_MPRJ[32] LA_DATA_IN_MPRJ[33] LA_DATA_IN_MPRJ[34] LA_DATA_IN_MPRJ[35] LA_DATA_IN_MPRJ[36] LA_DATA_IN_MPRJ[37] LA_DATA_IN_MPRJ[38] LA_DATA_IN_MPRJ[39] LA_DATA_IN_MPRJ[40] LA_DATA_IN_MPRJ[41] LA_DATA_IN_MPRJ[42] LA_DATA_IN_MPRJ[43] LA_DATA_IN_MPRJ[44] LA_DATA_IN_MPRJ[45] LA_DATA_IN_MPRJ[46] LA_DATA_IN_MPRJ[47] LA_DATA_IN_MPRJ[48] LA_DATA_IN_MPRJ[49] LA_DATA_IN_MPRJ[50] LA_DATA_IN_MPRJ[51] LA_DATA_IN_MPRJ[52] LA_DATA_IN_MPRJ[53] LA_DATA_IN_MPRJ[54] LA_DATA_IN_MPRJ[55] LA_DATA_IN_MPRJ[56] LA_DATA_IN_MPRJ[57] LA_DATA_IN_MPRJ[58] LA_DATA_IN_MPRJ[59] LA_DATA_IN_MPRJ[60] LA_DATA_IN_MPRJ[61] LA_DATA_IN_MPRJ[62] LA_DATA_IN_MPRJ[63] LA_DATA_IN_MPRJ[64] LA_DATA_IN_MPRJ[65] LA_DATA_IN_MPRJ[66] LA_DATA_IN_MPRJ[67] LA_DATA_IN_MPRJ[68] LA_DATA_IN_MPRJ[69] LA_DATA_IN_MPRJ[70] LA_DATA_IN_MPRJ[71] LA_DATA_IN_MPRJ[72] LA_DATA_IN_MPRJ[73] LA_DATA_IN_MPRJ[74] LA_DATA_IN_MPRJ[75] LA_DATA_IN_MPRJ[76] LA_DATA_IN_MPRJ[77] LA_DATA_IN_MPRJ[78] LA_DATA_IN_MPRJ[79] LA_DATA_IN_MPRJ[80] LA_DATA_IN_MPRJ[81] LA_DATA_IN_MPRJ[82] LA_DATA_IN_MPRJ[83] LA_DATA_IN_MPRJ[84] LA_DATA_IN_MPRJ[85] LA_DATA_IN_MPRJ[86] LA_DATA_IN_MPRJ[87] LA_DATA_IN_MPRJ[88] LA_DATA_IN_MPRJ[89] LA_DATA_IN_MPRJ[90] LA_DATA_IN_MPRJ[91] LA_DATA_IN_MPRJ[92] LA_DATA_IN_MPRJ[93] LA_DATA_IN_MPRJ[94] LA_DATA_IN_MPRJ[95] LA_DATA_IN_MPRJ[96] LA_DATA_IN_MPRJ[97] LA_DATA_IN_MPRJ[98] LA_DATA_IN_MPRJ[99] LA_DATA_IN_MPRJ[100] LA_DATA_IN_MPRJ[101] LA_DATA_IN_MPRJ[102] LA_DATA_IN_MPRJ[103] LA_DATA_IN_MPRJ[104] LA_DATA_IN_MPRJ[105] LA_DATA_IN_MPRJ[106] LA_DATA_IN_MPRJ[107] LA_DATA_IN_MPRJ[108] LA_DATA_IN_MPRJ[109] LA_DATA_IN_MPRJ[110] LA_DATA_IN_MPRJ[111] LA_DATA_IN_MPRJ[112] LA_DATA_IN_MPRJ[113] LA_DATA_IN_MPRJ[114] LA_DATA_IN_MPRJ[115] LA_DATA_IN_MPRJ[116] LA_DATA_IN_MPRJ[117] LA_DATA_IN_MPRJ[118] LA_DATA_IN_MPRJ[119] LA_DATA_IN_MPRJ[120] LA_DATA_IN_MPRJ[121] LA_DATA_IN_MPRJ[122] LA_DATA_IN_MPRJ[123] LA_DATA_IN_MPRJ[124] LA_DATA_IN_MPRJ[125] LA_DATA_IN_MPRJ[126] LA_DATA_IN_MPRJ[127] LA_DATA_OUT_CORE[0] LA_DATA_OUT_CORE[1] LA_DATA_OUT_CORE[2] LA_DATA_OUT_CORE[3] LA_DATA_OUT_CORE[4] LA_DATA_OUT_CORE[5] LA_DATA_OUT_CORE[6] LA_DATA_OUT_CORE[7] LA_DATA_OUT_CORE[8] LA_DATA_OUT_CORE[9] LA_DATA_OUT_CORE[10] LA_DATA_OUT_CORE[11] LA_DATA_OUT_CORE[12] LA_DATA_OUT_CORE[13] LA_DATA_OUT_CORE[14] LA_DATA_OUT_CORE[15] LA_DATA_OUT_CORE[16] LA_DATA_OUT_CORE[17] LA_DATA_OUT_CORE[18] LA_DATA_OUT_CORE[19] LA_DATA_OUT_CORE[20] LA_DATA_OUT_CORE[21] LA_DATA_OUT_CORE[22] LA_DATA_OUT_CORE[23] LA_DATA_OUT_CORE[24] LA_DATA_OUT_CORE[25] LA_DATA_OUT_CORE[26] LA_DATA_OUT_CORE[27] LA_DATA_OUT_CORE[28] LA_DATA_OUT_CORE[29] LA_DATA_OUT_CORE[30] LA_DATA_OUT_CORE[31] LA_DATA_OUT_CORE[32] LA_DATA_OUT_CORE[33] LA_DATA_OUT_CORE[34] LA_DATA_OUT_CORE[35] LA_DATA_OUT_CORE[36] LA_DATA_OUT_CORE[37] LA_DATA_OUT_CORE[38] LA_DATA_OUT_CORE[39] LA_DATA_OUT_CORE[40] LA_DATA_OUT_CORE[41] LA_DATA_OUT_CORE[42] LA_DATA_OUT_CORE[43] LA_DATA_OUT_CORE[44] LA_DATA_OUT_CORE[45] LA_DATA_OUT_CORE[46] LA_DATA_OUT_CORE[47] LA_DATA_OUT_CORE[48] LA_DATA_OUT_CORE[49] LA_DATA_OUT_CORE[50] LA_DATA_OUT_CORE[51] LA_DATA_OUT_CORE[52] LA_DATA_OUT_CORE[53] LA_DATA_OUT_CORE[54] LA_DATA_OUT_CORE[55] LA_DATA_OUT_CORE[56] LA_DATA_OUT_CORE[57] LA_DATA_OUT_CORE[58] LA_DATA_OUT_CORE[59] LA_DATA_OUT_CORE[60] LA_DATA_OUT_CORE[61] LA_DATA_OUT_CORE[62] LA_DATA_OUT_CORE[63] LA_DATA_OUT_CORE[64] LA_DATA_OUT_CORE[65] LA_DATA_OUT_CORE[66] LA_DATA_OUT_CORE[67] LA_DATA_OUT_CORE[68] LA_DATA_OUT_CORE[69] LA_DATA_OUT_CORE[70] LA_DATA_OUT_CORE[71] LA_DATA_OUT_CORE[72] LA_DATA_OUT_CORE[73] LA_DATA_OUT_CORE[74] LA_DATA_OUT_CORE[75] LA_DATA_OUT_CORE[76] LA_DATA_OUT_CORE[77] LA_DATA_OUT_CORE[78] LA_DATA_OUT_CORE[79] LA_DATA_OUT_CORE[80] LA_DATA_OUT_CORE[81] LA_DATA_OUT_CORE[82] LA_DATA_OUT_CORE[83] LA_DATA_OUT_CORE[84] LA_DATA_OUT_CORE[85] LA_DATA_OUT_CORE[86] LA_DATA_OUT_CORE[87] LA_DATA_OUT_CORE[88] LA_DATA_OUT_CORE[89] LA_DATA_OUT_CORE[90] LA_DATA_OUT_CORE[91] LA_DATA_OUT_CORE[92] LA_DATA_OUT_CORE[93] LA_DATA_OUT_CORE[94] LA_DATA_OUT_CORE[95] LA_DATA_OUT_CORE[96] LA_DATA_OUT_CORE[97] LA_DATA_OUT_CORE[98] LA_DATA_OUT_CORE[99] LA_DATA_OUT_CORE[100] LA_DATA_OUT_CORE[101] LA_DATA_OUT_CORE[102] LA_DATA_OUT_CORE[103] LA_DATA_OUT_CORE[104] LA_DATA_OUT_CORE[105] LA_DATA_OUT_CORE[106] LA_DATA_OUT_CORE[107] LA_DATA_OUT_CORE[108] LA_DATA_OUT_CORE[109] LA_DATA_OUT_CORE[110] LA_DATA_OUT_CORE[111] LA_DATA_OUT_CORE[112] LA_DATA_OUT_CORE[113] LA_DATA_OUT_CORE[114] LA_DATA_OUT_CORE[115] LA_DATA_OUT_CORE[116] LA_DATA_OUT_CORE[117] LA_DATA_OUT_CORE[118] LA_DATA_OUT_CORE[119] LA_DATA_OUT_CORE[120] LA_DATA_OUT_CORE[121] LA_DATA_OUT_CORE[122] LA_DATA_OUT_CORE[123] LA_DATA_OUT_CORE[124] LA_DATA_OUT_CORE[125] LA_DATA_OUT_CORE[126] LA_DATA_OUT_CORE[127] LA_DATA_OUT_MPRJ[0] LA_DATA_OUT_MPRJ[1] LA_DATA_OUT_MPRJ[2] LA_DATA_OUT_MPRJ[3] LA_DATA_OUT_MPRJ[4] LA_DATA_OUT_MPRJ[5] LA_DATA_OUT_MPRJ[6] LA_DATA_OUT_MPRJ[7] LA_DATA_OUT_MPRJ[8] LA_DATA_OUT_MPRJ[9] LA_DATA_OUT_MPRJ[10] LA_DATA_OUT_MPRJ[11] LA_DATA_OUT_MPRJ[12] LA_DATA_OUT_MPRJ[13] LA_DATA_OUT_MPRJ[14] LA_DATA_OUT_MPRJ[15] LA_DATA_OUT_MPRJ[16] LA_DATA_OUT_MPRJ[17] LA_DATA_OUT_MPRJ[18] LA_DATA_OUT_MPRJ[19] LA_DATA_OUT_MPRJ[20] LA_DATA_OUT_MPRJ[21] LA_DATA_OUT_MPRJ[22] LA_DATA_OUT_MPRJ[23] LA_DATA_OUT_MPRJ[24] LA_DATA_OUT_MPRJ[25] LA_DATA_OUT_MPRJ[26] LA_DATA_OUT_MPRJ[27] LA_DATA_OUT_MPRJ[28] LA_DATA_OUT_MPRJ[29] LA_DATA_OUT_MPRJ[30] LA_DATA_OUT_MPRJ[31] LA_DATA_OUT_MPRJ[32] LA_DATA_OUT_MPRJ[33] LA_DATA_OUT_MPRJ[34] LA_DATA_OUT_MPRJ[35] LA_DATA_OUT_MPRJ[36] LA_DATA_OUT_MPRJ[37] LA_DATA_OUT_MPRJ[38] LA_DATA_OUT_MPRJ[39] LA_DATA_OUT_MPRJ[40] LA_DATA_OUT_MPRJ[41] LA_DATA_OUT_MPRJ[42] LA_DATA_OUT_MPRJ[43] LA_DATA_OUT_MPRJ[44] LA_DATA_OUT_MPRJ[45] LA_DATA_OUT_MPRJ[46] LA_DATA_OUT_MPRJ[47] LA_DATA_OUT_MPRJ[48] LA_DATA_OUT_MPRJ[49] LA_DATA_OUT_MPRJ[50] LA_DATA_OUT_MPRJ[51] LA_DATA_OUT_MPRJ[52] LA_DATA_OUT_MPRJ[53] LA_DATA_OUT_MPRJ[54] LA_DATA_OUT_MPRJ[55] LA_DATA_OUT_MPRJ[56] LA_DATA_OUT_MPRJ[57] LA_DATA_OUT_MPRJ[58] LA_DATA_OUT_MPRJ[59] LA_DATA_OUT_MPRJ[60] LA_DATA_OUT_MPRJ[61] LA_DATA_OUT_MPRJ[62] LA_DATA_OUT_MPRJ[63] LA_DATA_OUT_MPRJ[64] LA_DATA_OUT_MPRJ[65] LA_DATA_OUT_MPRJ[66] LA_DATA_OUT_MPRJ[67] LA_DATA_OUT_MPRJ[68] LA_DATA_OUT_MPRJ[69] LA_DATA_OUT_MPRJ[70] LA_DATA_OUT_MPRJ[71] LA_DATA_OUT_MPRJ[72] LA_DATA_OUT_MPRJ[73] LA_DATA_OUT_MPRJ[74] LA_DATA_OUT_MPRJ[75] LA_DATA_OUT_MPRJ[76] LA_DATA_OUT_MPRJ[77] LA_DATA_OUT_MPRJ[78] LA_DATA_OUT_MPRJ[79] LA_DATA_OUT_MPRJ[80] LA_DATA_OUT_MPRJ[81] LA_DATA_OUT_MPRJ[82] LA_DATA_OUT_MPRJ[83] LA_DATA_OUT_MPRJ[84] LA_DATA_OUT_MPRJ[85] LA_DATA_OUT_MPRJ[86] LA_DATA_OUT_MPRJ[87] LA_DATA_OUT_MPRJ[88] LA_DATA_OUT_MPRJ[89] LA_DATA_OUT_MPRJ[90] LA_DATA_OUT_MPRJ[91] LA_DATA_OUT_MPRJ[92] LA_DATA_OUT_MPRJ[93] LA_DATA_OUT_MPRJ[94] LA_DATA_OUT_MPRJ[95] LA_DATA_OUT_MPRJ[96] LA_DATA_OUT_MPRJ[97] LA_DATA_OUT_MPRJ[98] LA_DATA_OUT_MPRJ[99] LA_DATA_OUT_MPRJ[100] LA_DATA_OUT_MPRJ[101] LA_DATA_OUT_MPRJ[102] LA_DATA_OUT_MPRJ[103] LA_DATA_OUT_MPRJ[104] LA_DATA_OUT_MPRJ[105] LA_DATA_OUT_MPRJ[106] LA_DATA_OUT_MPRJ[107] LA_DATA_OUT_MPRJ[108] LA_DATA_OUT_MPRJ[109] LA_DATA_OUT_MPRJ[110] LA_DATA_OUT_MPRJ[111] LA_DATA_OUT_MPRJ[112] LA_DATA_OUT_MPRJ[113] LA_DATA_OUT_MPRJ[114] LA_DATA_OUT_MPRJ[115] LA_DATA_OUT_MPRJ[116] LA_DATA_OUT_MPRJ[117] LA_DATA_OUT_MPRJ[118] LA_DATA_OUT_MPRJ[119] LA_DATA_OUT_MPRJ[120] LA_DATA_OUT_MPRJ[121] LA_DATA_OUT_MPRJ[122] LA_DATA_OUT_MPRJ[123] LA_DATA_OUT_MPRJ[124] LA_DATA_OUT_MPRJ[125] LA_DATA_OUT_MPRJ[126] LA_DATA_OUT_MPRJ[127] LA_IENA_MPRJ[0] LA_IENA_MPRJ[1] LA_IENA_MPRJ[2] LA_IENA_MPRJ[3] LA_IENA_MPRJ[4] LA_IENA_MPRJ[5] LA_IENA_MPRJ[6] LA_IENA_MPRJ[7] LA_IENA_MPRJ[8] LA_IENA_MPRJ[9] LA_IENA_MPRJ[10] LA_IENA_MPRJ[11] LA_IENA_MPRJ[12] LA_IENA_MPRJ[13] LA_IENA_MPRJ[14] LA_IENA_MPRJ[15] LA_IENA_MPRJ[16] LA_IENA_MPRJ[17] LA_IENA_MPRJ[18] LA_IENA_MPRJ[19] LA_IENA_MPRJ[20] LA_IENA_MPRJ[21] LA_IENA_MPRJ[22] LA_IENA_MPRJ[23] LA_IENA_MPRJ[24] LA_IENA_MPRJ[25] LA_IENA_MPRJ[26] LA_IENA_MPRJ[27] LA_IENA_MPRJ[28] LA_IENA_MPRJ[29] LA_IENA_MPRJ[30] LA_IENA_MPRJ[31] LA_IENA_MPRJ[32] LA_IENA_MPRJ[33] LA_IENA_MPRJ[34] LA_IENA_MPRJ[35] LA_IENA_MPRJ[36] LA_IENA_MPRJ[37] LA_IENA_MPRJ[38] LA_IENA_MPRJ[39] LA_IENA_MPRJ[40] LA_IENA_MPRJ[41] LA_IENA_MPRJ[42] LA_IENA_MPRJ[43] LA_IENA_MPRJ[44] LA_IENA_MPRJ[45] LA_IENA_MPRJ[46] LA_IENA_MPRJ[47] LA_IENA_MPRJ[48] LA_IENA_MPRJ[49] LA_IENA_MPRJ[50] LA_IENA_MPRJ[51] LA_IENA_MPRJ[52] LA_IENA_MPRJ[53] LA_IENA_MPRJ[54] LA_IENA_MPRJ[55] LA_IENA_MPRJ[56] LA_IENA_MPRJ[57] LA_IENA_MPRJ[58] LA_IENA_MPRJ[59] LA_IENA_MPRJ[60] LA_IENA_MPRJ[61] LA_IENA_MPRJ[62] LA_IENA_MPRJ[63] LA_IENA_MPRJ[64] LA_IENA_MPRJ[65] LA_IENA_MPRJ[66] LA_IENA_MPRJ[67] LA_IENA_MPRJ[68] LA_IENA_MPRJ[69] LA_IENA_MPRJ[70] LA_IENA_MPRJ[71] LA_IENA_MPRJ[72] LA_IENA_MPRJ[73] LA_IENA_MPRJ[74] LA_IENA_MPRJ[75] LA_IENA_MPRJ[76] LA_IENA_MPRJ[77] LA_IENA_MPRJ[78] LA_IENA_MPRJ[79] LA_IENA_MPRJ[80] LA_IENA_MPRJ[81] LA_IENA_MPRJ[82] LA_IENA_MPRJ[83] LA_IENA_MPRJ[84] LA_IENA_MPRJ[85] LA_IENA_MPRJ[86] LA_IENA_MPRJ[87] LA_IENA_MPRJ[88] LA_IENA_MPRJ[89] LA_IENA_MPRJ[90] LA_IENA_MPRJ[91] LA_IENA_MPRJ[92] LA_IENA_MPRJ[93] LA_IENA_MPRJ[94] LA_IENA_MPRJ[95] LA_IENA_MPRJ[96] LA_IENA_MPRJ[97] LA_IENA_MPRJ[98] LA_IENA_MPRJ[99] LA_IENA_MPRJ[100] LA_IENA_MPRJ[101] LA_IENA_MPRJ[102] LA_IENA_MPRJ[103] LA_IENA_MPRJ[104] LA_IENA_MPRJ[105] LA_IENA_MPRJ[106] LA_IENA_MPRJ[107] LA_IENA_MPRJ[108] LA_IENA_MPRJ[109] LA_IENA_MPRJ[110] LA_IENA_MPRJ[111] LA_IENA_MPRJ[112] LA_IENA_MPRJ[113] LA_IENA_MPRJ[114] LA_IENA_MPRJ[115] LA_IENA_MPRJ[116] LA_IENA_MPRJ[117] LA_IENA_MPRJ[118] LA_IENA_MPRJ[119] LA_IENA_MPRJ[120] LA_IENA_MPRJ[121] LA_IENA_MPRJ[122] LA_IENA_MPRJ[123] LA_IENA_MPRJ[124] LA_IENA_MPRJ[125] LA_IENA_MPRJ[126] LA_IENA_MPRJ[127] LA_OENB_CORE[0] LA_OENB_CORE[1] LA_OENB_CORE[2] LA_OENB_CORE[3] LA_OENB_CORE[4] LA_OENB_CORE[5] LA_OENB_CORE[6] LA_OENB_CORE[7] LA_OENB_CORE[8] LA_OENB_CORE[9] LA_OENB_CORE[10] LA_OENB_CORE[11] LA_OENB_CORE[12] LA_OENB_CORE[13] LA_OENB_CORE[14] LA_OENB_CORE[15] LA_OENB_CORE[16] LA_OENB_CORE[17] LA_OENB_CORE[18] LA_OENB_CORE[19] LA_OENB_CORE[20] LA_OENB_CORE[21] LA_OENB_CORE[22] LA_OENB_CORE[23] LA_OENB_CORE[24] LA_OENB_CORE[25] LA_OENB_CORE[26] LA_OENB_CORE[27] LA_OENB_CORE[28] LA_OENB_CORE[29] LA_OENB_CORE[30] LA_OENB_CORE[31] LA_OENB_CORE[32] LA_OENB_CORE[33] LA_OENB_CORE[34] LA_OENB_CORE[35] LA_OENB_CORE[36] LA_OENB_CORE[37] LA_OENB_CORE[38] LA_OENB_CORE[39] LA_OENB_CORE[40] LA_OENB_CORE[41] LA_OENB_CORE[42] LA_OENB_CORE[43] LA_OENB_CORE[44] LA_OENB_CORE[45] LA_OENB_CORE[46] LA_OENB_CORE[47] LA_OENB_CORE[48] LA_OENB_CORE[49] LA_OENB_CORE[50] LA_OENB_CORE[51] LA_OENB_CORE[52] LA_OENB_CORE[53] LA_OENB_CORE[54] LA_OENB_CORE[55] LA_OENB_CORE[56] LA_OENB_CORE[57] LA_OENB_CORE[58] LA_OENB_CORE[59] LA_OENB_CORE[60] LA_OENB_CORE[61] LA_OENB_CORE[62] LA_OENB_CORE[63] LA_OENB_CORE[64] LA_OENB_CORE[65] LA_OENB_CORE[66] LA_OENB_CORE[67] LA_OENB_CORE[68] LA_OENB_CORE[69] LA_OENB_CORE[70] LA_OENB_CORE[71] LA_OENB_CORE[72] LA_OENB_CORE[73] LA_OENB_CORE[74] LA_OENB_CORE[75] LA_OENB_CORE[76] LA_OENB_CORE[77] LA_OENB_CORE[78] LA_OENB_CORE[79] LA_OENB_CORE[80] LA_OENB_CORE[81] LA_OENB_CORE[82] LA_OENB_CORE[83] LA_OENB_CORE[84] LA_OENB_CORE[85] LA_OENB_CORE[86] LA_OENB_CORE[87] LA_OENB_CORE[88] LA_OENB_CORE[89] LA_OENB_CORE[90] LA_OENB_CORE[91] LA_OENB_CORE[92] LA_OENB_CORE[93] LA_OENB_CORE[94] LA_OENB_CORE[95] LA_OENB_CORE[96] LA_OENB_CORE[97] LA_OENB_CORE[98] LA_OENB_CORE[99] LA_OENB_CORE[100] LA_OENB_CORE[101] LA_OENB_CORE[102] LA_OENB_CORE[103] LA_OENB_CORE[104] LA_OENB_CORE[105] LA_OENB_CORE[106] LA_OENB_CORE[107] LA_OENB_CORE[108] LA_OENB_CORE[109] LA_OENB_CORE[110] LA_OENB_CORE[111] LA_OENB_CORE[112] LA_OENB_CORE[113] LA_OENB_CORE[114] LA_OENB_CORE[115] LA_OENB_CORE[116] LA_OENB_CORE[117] LA_OENB_CORE[118] LA_OENB_CORE[119] LA_OENB_CORE[120] LA_OENB_CORE[121] LA_OENB_CORE[122] LA_OENB_CORE[123] LA_OENB_CORE[124] LA_OENB_CORE[125] LA_OENB_CORE[126] LA_OENB_CORE[127] LA_OENB_MPRJ[0] LA_OENB_MPRJ[1] LA_OENB_MPRJ[2] LA_OENB_MPRJ[3] LA_OENB_MPRJ[4] LA_OENB_MPRJ[5] LA_OENB_MPRJ[6] LA_OENB_MPRJ[7] LA_OENB_MPRJ[8] LA_OENB_MPRJ[9] LA_OENB_MPRJ[10] LA_OENB_MPRJ[11] LA_OENB_MPRJ[12] LA_OENB_MPRJ[13] LA_OENB_MPRJ[14] LA_OENB_MPRJ[15] LA_OENB_MPRJ[16] LA_OENB_MPRJ[17] LA_OENB_MPRJ[18] LA_OENB_MPRJ[19] LA_OENB_MPRJ[20] LA_OENB_MPRJ[21] LA_OENB_MPRJ[22] LA_OENB_MPRJ[23] LA_OENB_MPRJ[24] LA_OENB_MPRJ[25] LA_OENB_MPRJ[26] LA_OENB_MPRJ[27] LA_OENB_MPRJ[28] LA_OENB_MPRJ[29] LA_OENB_MPRJ[30] LA_OENB_MPRJ[31] LA_OENB_MPRJ[32] LA_OENB_MPRJ[33] LA_OENB_MPRJ[34] LA_OENB_MPRJ[35] LA_OENB_MPRJ[36] LA_OENB_MPRJ[37] LA_OENB_MPRJ[38] LA_OENB_MPRJ[39] LA_OENB_MPRJ[40] LA_OENB_MPRJ[41] LA_OENB_MPRJ[42] LA_OENB_MPRJ[43] LA_OENB_MPRJ[44] LA_OENB_MPRJ[45] LA_OENB_MPRJ[46] LA_OENB_MPRJ[47] LA_OENB_MPRJ[48] LA_OENB_MPRJ[49] LA_OENB_MPRJ[50] LA_OENB_MPRJ[51] LA_OENB_MPRJ[52] LA_OENB_MPRJ[53] LA_OENB_MPRJ[54] LA_OENB_MPRJ[55] LA_OENB_MPRJ[56] LA_OENB_MPRJ[57] LA_OENB_MPRJ[58] LA_OENB_MPRJ[59] LA_OENB_MPRJ[60] LA_OENB_MPRJ[61] LA_OENB_MPRJ[62] LA_OENB_MPRJ[63] LA_OENB_MPRJ[64] LA_OENB_MPRJ[65] LA_OENB_MPRJ[66] LA_OENB_MPRJ[67] LA_OENB_MPRJ[68] LA_OENB_MPRJ[69] LA_OENB_MPRJ[70] LA_OENB_MPRJ[71] LA_OENB_MPRJ[72] LA_OENB_MPRJ[73] LA_OENB_MPRJ[74] LA_OENB_MPRJ[75] LA_OENB_MPRJ[76] LA_OENB_MPRJ[77] LA_OENB_MPRJ[78] LA_OENB_MPRJ[79] LA_OENB_MPRJ[80] LA_OENB_MPRJ[81] LA_OENB_MPRJ[82] LA_OENB_MPRJ[83] LA_OENB_MPRJ[84] LA_OENB_MPRJ[85] LA_OENB_MPRJ[86] LA_OENB_MPRJ[87] LA_OENB_MPRJ[88] LA_OENB_MPRJ[89] LA_OENB_MPRJ[90] LA_OENB_MPRJ[91] LA_OENB_MPRJ[92] LA_OENB_MPRJ[93] LA_OENB_MPRJ[94] LA_OENB_MPRJ[95] LA_OENB_MPRJ[96] LA_OENB_MPRJ[97] LA_OENB_MPRJ[98] LA_OENB_MPRJ[99] LA_OENB_MPRJ[100] LA_OENB_MPRJ[101] LA_OENB_MPRJ[102] LA_OENB_MPRJ[103] LA_OENB_MPRJ[104] LA_OENB_MPRJ[105] LA_OENB_MPRJ[106] LA_OENB_MPRJ[107] LA_OENB_MPRJ[108] LA_OENB_MPRJ[109] LA_OENB_MPRJ[110] LA_OENB_MPRJ[111] LA_OENB_MPRJ[112] LA_OENB_MPRJ[113] LA_OENB_MPRJ[114] LA_OENB_MPRJ[115] LA_OENB_MPRJ[116] LA_OENB_MPRJ[117] LA_OENB_MPRJ[118] LA_OENB_MPRJ[119] LA_OENB_MPRJ[120] LA_OENB_MPRJ[121] LA_OENB_MPRJ[122] LA_OENB_MPRJ[123] LA_OENB_MPRJ[124] LA_OENB_MPRJ[125] LA_OENB_MPRJ[126] LA_OENB_MPRJ[127] MPRJ_ADR_O_CORE[0] MPRJ_ADR_O_CORE[1] MPRJ_ADR_O_CORE[2] MPRJ_ADR_O_CORE[3] MPRJ_ADR_O_CORE[4] MPRJ_ADR_O_CORE[5] MPRJ_ADR_O_CORE[6] MPRJ_ADR_O_CORE[7] MPRJ_ADR_O_CORE[8] MPRJ_ADR_O_CORE[9] MPRJ_ADR_O_CORE[10] MPRJ_ADR_O_CORE[11] MPRJ_ADR_O_CORE[12] MPRJ_ADR_O_CORE[13] MPRJ_ADR_O_CORE[14] MPRJ_ADR_O_CORE[15] MPRJ_ADR_O_CORE[16] MPRJ_ADR_O_CORE[17] MPRJ_ADR_O_CORE[18] MPRJ_ADR_O_CORE[19] MPRJ_ADR_O_CORE[20] MPRJ_ADR_O_CORE[21] MPRJ_ADR_O_CORE[22] MPRJ_ADR_O_CORE[23] MPRJ_ADR_O_CORE[24] MPRJ_ADR_O_CORE[25] MPRJ_ADR_O_CORE[26] MPRJ_ADR_O_CORE[27] MPRJ_ADR_O_CORE[28] MPRJ_ADR_O_CORE[29] MPRJ_ADR_O_CORE[30] MPRJ_ADR_O_CORE[31] MPRJ_ADR_O_USER[0] MPRJ_ADR_O_USER[1] MPRJ_ADR_O_USER[2] MPRJ_ADR_O_USER[3] MPRJ_ADR_O_USER[4] MPRJ_ADR_O_USER[5] MPRJ_ADR_O_USER[6] MPRJ_ADR_O_USER[7] MPRJ_ADR_O_USER[8] MPRJ_ADR_O_USER[9] MPRJ_ADR_O_USER[10] MPRJ_ADR_O_USER[11] MPRJ_ADR_O_USER[12] MPRJ_ADR_O_USER[13] MPRJ_ADR_O_USER[14] MPRJ_ADR_O_USER[15] MPRJ_ADR_O_USER[16] MPRJ_ADR_O_USER[17] MPRJ_ADR_O_USER[18] MPRJ_ADR_O_USER[19] MPRJ_ADR_O_USER[20] MPRJ_ADR_O_USER[21] MPRJ_ADR_O_USER[22] MPRJ_ADR_O_USER[23] MPRJ_ADR_O_USER[24] MPRJ_ADR_O_USER[25] MPRJ_ADR_O_USER[26] MPRJ_ADR_O_USER[27] MPRJ_ADR_O_USER[28] MPRJ_ADR_O_USER[29] MPRJ_ADR_O_USER[30] MPRJ_ADR_O_USER[31] MPRJ_DAT_I_CORE[0] MPRJ_DAT_I_CORE[1] MPRJ_DAT_I_CORE[2] MPRJ_DAT_I_CORE[3] MPRJ_DAT_I_CORE[4] MPRJ_DAT_I_CORE[5] MPRJ_DAT_I_CORE[6] MPRJ_DAT_I_CORE[7] MPRJ_DAT_I_CORE[8] MPRJ_DAT_I_CORE[9] MPRJ_DAT_I_CORE[10] MPRJ_DAT_I_CORE[11] MPRJ_DAT_I_CORE[12] MPRJ_DAT_I_CORE[13] MPRJ_DAT_I_CORE[14] MPRJ_DAT_I_CORE[15] MPRJ_DAT_I_CORE[16] MPRJ_DAT_I_CORE[17] MPRJ_DAT_I_CORE[18] MPRJ_DAT_I_CORE[19] MPRJ_DAT_I_CORE[20] MPRJ_DAT_I_CORE[21] MPRJ_DAT_I_CORE[22] MPRJ_DAT_I_CORE[23] MPRJ_DAT_I_CORE[24] MPRJ_DAT_I_CORE[25] MPRJ_DAT_I_CORE[26] MPRJ_DAT_I_CORE[27] MPRJ_DAT_I_CORE[28] MPRJ_DAT_I_CORE[29] MPRJ_DAT_I_CORE[30] MPRJ_DAT_I_CORE[31] MPRJ_DAT_I_USER[0] MPRJ_DAT_I_USER[1] MPRJ_DAT_I_USER[2] MPRJ_DAT_I_USER[3] MPRJ_DAT_I_USER[4] MPRJ_DAT_I_USER[5] MPRJ_DAT_I_USER[6] MPRJ_DAT_I_USER[7] MPRJ_DAT_I_USER[8] MPRJ_DAT_I_USER[9] MPRJ_DAT_I_USER[10] MPRJ_DAT_I_USER[11] MPRJ_DAT_I_USER[12] MPRJ_DAT_I_USER[13] MPRJ_DAT_I_USER[14] MPRJ_DAT_I_USER[15] MPRJ_DAT_I_USER[16] MPRJ_DAT_I_USER[17] MPRJ_DAT_I_USER[18] MPRJ_DAT_I_USER[19] MPRJ_DAT_I_USER[20] MPRJ_DAT_I_USER[21] MPRJ_DAT_I_USER[22] MPRJ_DAT_I_USER[23] MPRJ_DAT_I_USER[24] MPRJ_DAT_I_USER[25] MPRJ_DAT_I_USER[26] MPRJ_DAT_I_USER[27] MPRJ_DAT_I_USER[28] MPRJ_DAT_I_USER[29] MPRJ_DAT_I_USER[30] MPRJ_DAT_I_USER[31] MPRJ_DAT_O_CORE[0] MPRJ_DAT_O_CORE[1] MPRJ_DAT_O_CORE[2] MPRJ_DAT_O_CORE[3] MPRJ_DAT_O_CORE[4] MPRJ_DAT_O_CORE[5] MPRJ_DAT_O_CORE[6] MPRJ_DAT_O_CORE[7] MPRJ_DAT_O_CORE[8] MPRJ_DAT_O_CORE[9] MPRJ_DAT_O_CORE[10] MPRJ_DAT_O_CORE[11] MPRJ_DAT_O_CORE[12] MPRJ_DAT_O_CORE[13] MPRJ_DAT_O_CORE[14] MPRJ_DAT_O_CORE[15] MPRJ_DAT_O_CORE[16] MPRJ_DAT_O_CORE[17] MPRJ_DAT_O_CORE[18] MPRJ_DAT_O_CORE[19] MPRJ_DAT_O_CORE[20] MPRJ_DAT_O_CORE[21] MPRJ_DAT_O_CORE[22] MPRJ_DAT_O_CORE[23] MPRJ_DAT_O_CORE[24] MPRJ_DAT_O_CORE[25] MPRJ_DAT_O_CORE[26] MPRJ_DAT_O_CORE[27] MPRJ_DAT_O_CORE[28] MPRJ_DAT_O_CORE[29] MPRJ_DAT_O_CORE[30] MPRJ_DAT_O_CORE[31] MPRJ_DAT_O_USER[0] MPRJ_DAT_O_USER[1] MPRJ_DAT_O_USER[2] MPRJ_DAT_O_USER[3] MPRJ_DAT_O_USER[4] MPRJ_DAT_O_USER[5] MPRJ_DAT_O_USER[6] MPRJ_DAT_O_USER[7] MPRJ_DAT_O_USER[8] MPRJ_DAT_O_USER[9] MPRJ_DAT_O_USER[10] MPRJ_DAT_O_USER[11] MPRJ_DAT_O_USER[12] MPRJ_DAT_O_USER[13] MPRJ_DAT_O_USER[14] MPRJ_DAT_O_USER[15] MPRJ_DAT_O_USER[16] MPRJ_DAT_O_USER[17] MPRJ_DAT_O_USER[18] MPRJ_DAT_O_USER[19] MPRJ_DAT_O_USER[20] MPRJ_DAT_O_USER[21] MPRJ_DAT_O_USER[22] MPRJ_DAT_O_USER[23] MPRJ_DAT_O_USER[24] MPRJ_DAT_O_USER[25] MPRJ_DAT_O_USER[26] MPRJ_DAT_O_USER[27] MPRJ_DAT_O_USER[28] MPRJ_DAT_O_USER[29] MPRJ_DAT_O_USER[30] MPRJ_DAT_O_USER[31] MPRJ_SEL_O_CORE[0] MPRJ_SEL_O_CORE[1] MPRJ_SEL_O_CORE[2] MPRJ_SEL_O_CORE[3] MPRJ_SEL_O_USER[0] MPRJ_SEL_O_USER[1] MPRJ_SEL_O_USER[2] MPRJ_SEL_O_USER[3] USER_IRQ[0] USER_IRQ[1] USER_IRQ[2] USER_IRQ_CORE[0] USER_IRQ_CORE[1] USER_IRQ_CORE[2] USER_IRQ_ENA[0] USER_IRQ_ENA[1] USER_IRQ_ENA[2] 

XANTENNA__329__A NET478 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__330__A NET479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__331__A NET480 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__332__A NET481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__333__A NET483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__334__A NET484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__335__A NET485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__336__A NET486 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__337__A NET487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__338__A NET488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__339__A NET489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__340__A NET490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__341__A NET491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__342__A NET492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__343__A NET494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__344__A NET495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__345__A NET496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__346__A NET497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__347__A NET498 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__348__A NET499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__349__A NET500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__350__A NET501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__351__A NET502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__352__A NET503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__353__A NET505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__354__A NET506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__355__A NET507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__356__A NET508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__357__A NET509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__358__A NET510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__359__A NET511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__360__A NET512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__361__A NET513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__362__A NET514 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__363__A NET389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__364__A NET390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__365__A NET391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__366__A NET392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__367__A NET393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__368__A NET394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__369__A NET395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__370__A NET396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__371__A NET397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__372__A NET398 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__373__A NET400 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__374__A NET401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__375__A NET402 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__376__A NET403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__377__A NET404 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__378__A NET405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__379__A NET406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__380__A NET407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__381__A NET408 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__382__A NET409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__383__A NET411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__384__A NET412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__385__A NET413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__386__A NET414 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__387__A NET415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__388__A NET416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__389__A NET417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__390__A NET418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__391__A NET1 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__392__A NET2 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__393__A NET549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__394__A NET619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__395__A NET620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__396__A NET615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__397__A NET616 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__398__A NET617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__399__A NET618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__400__A NET517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__401__A NET528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__402__A NET539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__403__A NET542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__404__A NET543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__405__A NET544 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__406__A NET545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__407__A NET546 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__408__A NET547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__409__A NET548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__410__A NET518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__411__A NET519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__412__A NET520 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__413__A NET521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__414__A NET522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__415__A NET523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__416__A NET524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__417__A NET525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__418__A NET526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__419__A NET527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__420__A NET529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__421__A NET530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__422__A NET531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__423__A NET532 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__424__A NET533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__425__A NET534 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__426__A NET535 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__427__A NET536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__428__A NET537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__429__A NET538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__430__A NET540 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__431__A NET541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__432__A NET582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__433__A NET593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__434__A NET604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__435__A NET607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__436__A NET608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__437__A NET609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__438__A NET610 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__439__A NET611 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__440__A NET612 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__441__A NET613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__442__A NET583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__443__A NET584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__444__A NET585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__445__A NET586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__446__A NET587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__447__A NET588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__448__A NET589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__449__A NET590 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__450__A NET591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__451__A NET592 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__452__A NET594 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__453__A NET595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__454__A NET596 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__455__A NET597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__456__A NET598 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__457__A NET599 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__458__A NET600 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__459__A NET601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__460__A NET602 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__461__A NET603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__462__A NET605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__463__A NET606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__464__A NET132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__465__A NET171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__466__A NET182 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__467__A NET193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__468__A NET204 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__469__A NET215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__470__A NET226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__471__A NET237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__472__A NET248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__473__A NET259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__474__A NET143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__475__A NET154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__476__A NET163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__477__A NET164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__478__A NET165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__479__A NET166 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__480__A NET167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__481__A NET168 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__482__A NET169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__483__A NET170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__484__A NET172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__485__A NET173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__486__A NET174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__487__A NET175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__488__A NET176 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__489__A NET177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__490__A NET178 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__491__A NET179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__492__A NET180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__493__A NET181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__494__A NET183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__495__A NET184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__496__A NET185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__497__A NET186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__498__A NET187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__499__A NET188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__500__A NET189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__501__A NET190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__502__A NET191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__503__A NET192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__504__A NET194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__505__A NET195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__506__A NET196 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__507__A NET197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__508__A NET198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__509__A NET199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__510__A NET200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__511__A NET201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__512__A NET202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__513__A NET203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__514__A NET205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__515__A NET206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__516__A NET207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__517__A NET208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__518__A NET209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__519__A NET210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__520__A NET211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__521__A NET212 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__522__A NET213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__523__A NET214 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__524__A NET216 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__525__A NET217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__526__A NET218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__527__A NET219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__528__A NET220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__529__A NET221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__530__A NET222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__531__A NET223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__532__A NET224 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__533__A NET225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__534__A NET227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__535__A NET228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__536__A NET229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__537__A NET230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__538__A NET231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__539__A NET232 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__540__A NET233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__541__A NET234 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__542__A NET235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__543__A NET236 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__544__A NET238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__545__A NET239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__546__A NET240 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__547__A NET241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__548__A NET242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__549__A NET243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__550__A NET244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__551__A NET245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__552__A NET246 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__553__A NET247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__554__A NET249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__555__A NET250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__556__A NET251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__557__A NET252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__558__A NET253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__559__A NET254 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__560__A NET255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__561__A NET256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__562__A NET257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__563__A NET258 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__564__A NET133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__565__A NET134 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__566__A NET135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__567__A NET136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__568__A NET137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__569__A NET138 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__570__A NET139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__571__A NET140 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__572__A NET141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__573__A NET142 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__574__A NET144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__575__A NET145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__576__A NET146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__577__A NET147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__578__A NET148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__579__A NET149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__580__A NET150 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__581__A NET151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__582__A NET152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__583__A NET153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__584__A NET155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__585__A NET156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__586__A NET157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__587__A NET158 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__588__A NET159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__589__A NET160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__590__A NET161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__591__A NET162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__592__A NET388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__593__A NET427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__594__A NET438 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__595__A NET449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__596__A NET460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__597__A NET471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__598__A NET482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__599__A NET493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__600__A NET504 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__601__A NET515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__602__A NET399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__603__A NET410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__604__A NET419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__605__A NET420 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__606__A NET421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__607__A NET422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__608__A NET423 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__609__A NET424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__610__A NET425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__611__A NET426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__612__A NET428 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__613__A NET429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__614__A NET430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__615__A NET431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__616__A NET432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__617__A NET433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__618__A NET434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__619__A NET435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__620__A NET436 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__621__A NET437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__622__A NET439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__623__A NET440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__624__A NET441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__625__A NET442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__626__A NET443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__627__A NET444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__628__A NET445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__629__A NET446 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__630__A NET447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__631__A NET448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__632__A NET450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__633__A NET451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__634__A NET452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__635__A NET453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__636__A NET454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__637__A NET455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__638__A NET456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__639__A NET457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__640__A NET458 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__641__A NET459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__642__A NET461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__643__A NET462 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__644__A NET463 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__645__A NET464 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__646__A NET465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__647__A NET466 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__648__A NET467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__649__A NET468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__650__A NET469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__651__A NET470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__652__A NET472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__653__A NET473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__654__A NET474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__655__A NET475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__656__A NET476 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA__657__A NET477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT100_A LA_DATA_OUT_CORE[71] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT101_A LA_DATA_OUT_CORE[72] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT102_A LA_DATA_OUT_CORE[73] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT103_A LA_DATA_OUT_CORE[74] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT104_A LA_DATA_OUT_CORE[75] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT105_A LA_DATA_OUT_CORE[76] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT106_A LA_DATA_OUT_CORE[77] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT107_A LA_DATA_OUT_CORE[78] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT108_A LA_DATA_OUT_CORE[79] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT109_A LA_DATA_OUT_CORE[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT10_A LA_DATA_OUT_CORE[105] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT110_A LA_DATA_OUT_CORE[80] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT111_A LA_DATA_OUT_CORE[81] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT112_A LA_DATA_OUT_CORE[82] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT113_A LA_DATA_OUT_CORE[83] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT114_A LA_DATA_OUT_CORE[84] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT115_A LA_DATA_OUT_CORE[85] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT116_A LA_DATA_OUT_CORE[86] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT117_A LA_DATA_OUT_CORE[87] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT118_A LA_DATA_OUT_CORE[88] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT119_A LA_DATA_OUT_CORE[89] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT11_A LA_DATA_OUT_CORE[106] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT120_A LA_DATA_OUT_CORE[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT121_A LA_DATA_OUT_CORE[90] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT122_A LA_DATA_OUT_CORE[91] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT123_A LA_DATA_OUT_CORE[92] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT124_A LA_DATA_OUT_CORE[93] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT125_A LA_DATA_OUT_CORE[94] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT126_A LA_DATA_OUT_CORE[95] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT127_A LA_DATA_OUT_CORE[96] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT128_A LA_DATA_OUT_CORE[97] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT129_A LA_DATA_OUT_CORE[98] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT12_A LA_DATA_OUT_CORE[107] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT130_A LA_DATA_OUT_CORE[99] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT131_A LA_DATA_OUT_CORE[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT132_A LA_DATA_OUT_MPRJ[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT133_A LA_DATA_OUT_MPRJ[100] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT134_A LA_DATA_OUT_MPRJ[101] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT135_A LA_DATA_OUT_MPRJ[102] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT136_A LA_DATA_OUT_MPRJ[103] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT137_A LA_DATA_OUT_MPRJ[104] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT138_A LA_DATA_OUT_MPRJ[105] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT139_A LA_DATA_OUT_MPRJ[106] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT13_A LA_DATA_OUT_CORE[108] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT140_A LA_DATA_OUT_MPRJ[107] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT141_A LA_DATA_OUT_MPRJ[108] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT142_A LA_DATA_OUT_MPRJ[109] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT143_A LA_DATA_OUT_MPRJ[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT144_A LA_DATA_OUT_MPRJ[110] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT145_A LA_DATA_OUT_MPRJ[111] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT146_A LA_DATA_OUT_MPRJ[112] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT147_A LA_DATA_OUT_MPRJ[113] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT148_A LA_DATA_OUT_MPRJ[114] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT149_A LA_DATA_OUT_MPRJ[115] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT14_A LA_DATA_OUT_CORE[109] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT150_A LA_DATA_OUT_MPRJ[116] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT151_A LA_DATA_OUT_MPRJ[117] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT152_A LA_DATA_OUT_MPRJ[118] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT153_A LA_DATA_OUT_MPRJ[119] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT154_A LA_DATA_OUT_MPRJ[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT155_A LA_DATA_OUT_MPRJ[120] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT156_A LA_DATA_OUT_MPRJ[121] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT157_A LA_DATA_OUT_MPRJ[122] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT158_A LA_DATA_OUT_MPRJ[123] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT159_A LA_DATA_OUT_MPRJ[124] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT15_A LA_DATA_OUT_CORE[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT160_A LA_DATA_OUT_MPRJ[125] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT161_A LA_DATA_OUT_MPRJ[126] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT162_A LA_DATA_OUT_MPRJ[127] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT163_A LA_DATA_OUT_MPRJ[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT164_A LA_DATA_OUT_MPRJ[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT165_A LA_DATA_OUT_MPRJ[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT166_A LA_DATA_OUT_MPRJ[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT167_A LA_DATA_OUT_MPRJ[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT168_A LA_DATA_OUT_MPRJ[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT169_A LA_DATA_OUT_MPRJ[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT16_A LA_DATA_OUT_CORE[110] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT170_A LA_DATA_OUT_MPRJ[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT171_A LA_DATA_OUT_MPRJ[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT172_A LA_DATA_OUT_MPRJ[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT173_A LA_DATA_OUT_MPRJ[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT174_A LA_DATA_OUT_MPRJ[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT175_A LA_DATA_OUT_MPRJ[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT176_A LA_DATA_OUT_MPRJ[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT177_A LA_DATA_OUT_MPRJ[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT178_A LA_DATA_OUT_MPRJ[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT179_A LA_DATA_OUT_MPRJ[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT17_A LA_DATA_OUT_CORE[111] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT180_A LA_DATA_OUT_MPRJ[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT181_A LA_DATA_OUT_MPRJ[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT182_A LA_DATA_OUT_MPRJ[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT183_A LA_DATA_OUT_MPRJ[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT184_A LA_DATA_OUT_MPRJ[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT185_A LA_DATA_OUT_MPRJ[32] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT186_A LA_DATA_OUT_MPRJ[33] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT187_A LA_DATA_OUT_MPRJ[34] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT188_A LA_DATA_OUT_MPRJ[35] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT189_A LA_DATA_OUT_MPRJ[36] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT18_A LA_DATA_OUT_CORE[112] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT190_A LA_DATA_OUT_MPRJ[37] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT191_A LA_DATA_OUT_MPRJ[38] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT192_A LA_DATA_OUT_MPRJ[39] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT193_A LA_DATA_OUT_MPRJ[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT194_A LA_DATA_OUT_MPRJ[40] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT195_A LA_DATA_OUT_MPRJ[41] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT196_A LA_DATA_OUT_MPRJ[42] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT197_A LA_DATA_OUT_MPRJ[43] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT198_A LA_DATA_OUT_MPRJ[44] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT199_A LA_DATA_OUT_MPRJ[45] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT19_A LA_DATA_OUT_CORE[113] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT1_A CARAVEL_CLK VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT200_A LA_DATA_OUT_MPRJ[46] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT201_A LA_DATA_OUT_MPRJ[47] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT202_A LA_DATA_OUT_MPRJ[48] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT203_A LA_DATA_OUT_MPRJ[49] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT204_A LA_DATA_OUT_MPRJ[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT205_A LA_DATA_OUT_MPRJ[50] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT206_A LA_DATA_OUT_MPRJ[51] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT207_A LA_DATA_OUT_MPRJ[52] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT208_A LA_DATA_OUT_MPRJ[53] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT209_A LA_DATA_OUT_MPRJ[54] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT20_A LA_DATA_OUT_CORE[114] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT210_A LA_DATA_OUT_MPRJ[55] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT211_A LA_DATA_OUT_MPRJ[56] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT212_A LA_DATA_OUT_MPRJ[57] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT213_A LA_DATA_OUT_MPRJ[58] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT214_A LA_DATA_OUT_MPRJ[59] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT215_A LA_DATA_OUT_MPRJ[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT216_A LA_DATA_OUT_MPRJ[60] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT217_A LA_DATA_OUT_MPRJ[61] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT218_A LA_DATA_OUT_MPRJ[62] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT219_A LA_DATA_OUT_MPRJ[63] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT21_A LA_DATA_OUT_CORE[115] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT220_A LA_DATA_OUT_MPRJ[64] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT221_A LA_DATA_OUT_MPRJ[65] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT222_A LA_DATA_OUT_MPRJ[66] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT223_A LA_DATA_OUT_MPRJ[67] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT224_A LA_DATA_OUT_MPRJ[68] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT225_A LA_DATA_OUT_MPRJ[69] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT226_A LA_DATA_OUT_MPRJ[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT227_A LA_DATA_OUT_MPRJ[70] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT228_A LA_DATA_OUT_MPRJ[71] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT229_A LA_DATA_OUT_MPRJ[72] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT22_A LA_DATA_OUT_CORE[116] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT230_A LA_DATA_OUT_MPRJ[73] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT231_A LA_DATA_OUT_MPRJ[74] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT232_A LA_DATA_OUT_MPRJ[75] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT233_A LA_DATA_OUT_MPRJ[76] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT234_A LA_DATA_OUT_MPRJ[77] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT235_A LA_DATA_OUT_MPRJ[78] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT236_A LA_DATA_OUT_MPRJ[79] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT237_A LA_DATA_OUT_MPRJ[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT238_A LA_DATA_OUT_MPRJ[80] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT239_A LA_DATA_OUT_MPRJ[81] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT23_A LA_DATA_OUT_CORE[117] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT240_A LA_DATA_OUT_MPRJ[82] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT241_A LA_DATA_OUT_MPRJ[83] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT242_A LA_DATA_OUT_MPRJ[84] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT243_A LA_DATA_OUT_MPRJ[85] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT244_A LA_DATA_OUT_MPRJ[86] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT245_A LA_DATA_OUT_MPRJ[87] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT246_A LA_DATA_OUT_MPRJ[88] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT247_A LA_DATA_OUT_MPRJ[89] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT248_A LA_DATA_OUT_MPRJ[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT249_A LA_DATA_OUT_MPRJ[90] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT24_A LA_DATA_OUT_CORE[118] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT250_A LA_DATA_OUT_MPRJ[91] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT251_A LA_DATA_OUT_MPRJ[92] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT252_A LA_DATA_OUT_MPRJ[93] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT253_A LA_DATA_OUT_MPRJ[94] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT254_A LA_DATA_OUT_MPRJ[95] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT255_A LA_DATA_OUT_MPRJ[96] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT256_A LA_DATA_OUT_MPRJ[97] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT257_A LA_DATA_OUT_MPRJ[98] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT258_A LA_DATA_OUT_MPRJ[99] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT259_A LA_DATA_OUT_MPRJ[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT25_A LA_DATA_OUT_CORE[119] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT260_A LA_IENA_MPRJ[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT261_A LA_IENA_MPRJ[100] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT262_A LA_IENA_MPRJ[101] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT263_A LA_IENA_MPRJ[102] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT264_A LA_IENA_MPRJ[103] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT265_A LA_IENA_MPRJ[104] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT266_A LA_IENA_MPRJ[105] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT267_A LA_IENA_MPRJ[106] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT268_A LA_IENA_MPRJ[107] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT269_A LA_IENA_MPRJ[108] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT26_A LA_DATA_OUT_CORE[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT270_A LA_IENA_MPRJ[109] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT271_A LA_IENA_MPRJ[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT272_A LA_IENA_MPRJ[110] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT273_A LA_IENA_MPRJ[111] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT274_A LA_IENA_MPRJ[112] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT275_A LA_IENA_MPRJ[113] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT276_A LA_IENA_MPRJ[114] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT277_A LA_IENA_MPRJ[115] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT278_A LA_IENA_MPRJ[116] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT279_A LA_IENA_MPRJ[117] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT27_A LA_DATA_OUT_CORE[120] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT280_A LA_IENA_MPRJ[118] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT281_A LA_IENA_MPRJ[119] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT282_A LA_IENA_MPRJ[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT283_A LA_IENA_MPRJ[120] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT284_A LA_IENA_MPRJ[121] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT285_A LA_IENA_MPRJ[122] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT286_A LA_IENA_MPRJ[123] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT287_A LA_IENA_MPRJ[124] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT288_A LA_IENA_MPRJ[125] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT289_A LA_IENA_MPRJ[126] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT28_A LA_DATA_OUT_CORE[121] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT290_A LA_IENA_MPRJ[127] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT291_A LA_IENA_MPRJ[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT292_A LA_IENA_MPRJ[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT293_A LA_IENA_MPRJ[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT294_A LA_IENA_MPRJ[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT295_A LA_IENA_MPRJ[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT296_A LA_IENA_MPRJ[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT297_A LA_IENA_MPRJ[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT298_A LA_IENA_MPRJ[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT299_A LA_IENA_MPRJ[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT29_A LA_DATA_OUT_CORE[122] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT2_A CARAVEL_CLK2 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT300_A LA_IENA_MPRJ[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT301_A LA_IENA_MPRJ[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT302_A LA_IENA_MPRJ[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT303_A LA_IENA_MPRJ[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT304_A LA_IENA_MPRJ[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT305_A LA_IENA_MPRJ[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT306_A LA_IENA_MPRJ[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT307_A LA_IENA_MPRJ[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT308_A LA_IENA_MPRJ[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT309_A LA_IENA_MPRJ[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT30_A LA_DATA_OUT_CORE[123] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT310_A LA_IENA_MPRJ[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT311_A LA_IENA_MPRJ[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT312_A LA_IENA_MPRJ[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT313_A LA_IENA_MPRJ[32] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT314_A LA_IENA_MPRJ[33] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT315_A LA_IENA_MPRJ[34] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT316_A LA_IENA_MPRJ[35] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT317_A LA_IENA_MPRJ[36] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT318_A LA_IENA_MPRJ[37] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT319_A LA_IENA_MPRJ[38] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT31_A LA_DATA_OUT_CORE[124] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT320_A LA_IENA_MPRJ[39] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT321_A LA_IENA_MPRJ[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT322_A LA_IENA_MPRJ[40] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT323_A LA_IENA_MPRJ[41] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT324_A LA_IENA_MPRJ[42] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT325_A LA_IENA_MPRJ[43] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT326_A LA_IENA_MPRJ[44] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT327_A LA_IENA_MPRJ[45] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT328_A LA_IENA_MPRJ[46] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT329_A LA_IENA_MPRJ[47] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT32_A LA_DATA_OUT_CORE[125] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT330_A LA_IENA_MPRJ[48] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT331_A LA_IENA_MPRJ[49] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT332_A LA_IENA_MPRJ[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT333_A LA_IENA_MPRJ[50] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT334_A LA_IENA_MPRJ[51] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT335_A LA_IENA_MPRJ[52] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT336_A LA_IENA_MPRJ[53] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT337_A LA_IENA_MPRJ[54] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT338_A LA_IENA_MPRJ[55] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT339_A LA_IENA_MPRJ[56] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT33_A LA_DATA_OUT_CORE[126] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT340_A LA_IENA_MPRJ[57] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT341_A LA_IENA_MPRJ[58] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT342_A LA_IENA_MPRJ[59] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT343_A LA_IENA_MPRJ[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT344_A LA_IENA_MPRJ[60] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT345_A LA_IENA_MPRJ[61] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT346_A LA_IENA_MPRJ[62] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT347_A LA_IENA_MPRJ[63] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT348_A LA_IENA_MPRJ[64] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT349_A LA_IENA_MPRJ[65] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT34_A LA_DATA_OUT_CORE[127] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT350_A LA_IENA_MPRJ[66] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT351_A LA_IENA_MPRJ[67] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT352_A LA_IENA_MPRJ[68] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT353_A LA_IENA_MPRJ[69] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT354_A LA_IENA_MPRJ[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT355_A LA_IENA_MPRJ[70] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT356_A LA_IENA_MPRJ[71] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT357_A LA_IENA_MPRJ[72] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT358_A LA_IENA_MPRJ[73] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT359_A LA_IENA_MPRJ[74] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT35_A LA_DATA_OUT_CORE[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT360_A LA_IENA_MPRJ[75] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT361_A LA_IENA_MPRJ[76] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT362_A LA_IENA_MPRJ[77] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT363_A LA_IENA_MPRJ[78] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT364_A LA_IENA_MPRJ[79] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT365_A LA_IENA_MPRJ[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT366_A LA_IENA_MPRJ[80] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT367_A LA_IENA_MPRJ[81] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT368_A LA_IENA_MPRJ[82] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT369_A LA_IENA_MPRJ[83] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT36_A LA_DATA_OUT_CORE[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT370_A LA_IENA_MPRJ[84] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT371_A LA_IENA_MPRJ[85] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT372_A LA_IENA_MPRJ[86] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT373_A LA_IENA_MPRJ[87] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT374_A LA_IENA_MPRJ[88] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT375_A LA_IENA_MPRJ[89] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT376_A LA_IENA_MPRJ[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT377_A LA_IENA_MPRJ[90] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT378_A LA_IENA_MPRJ[91] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT379_A LA_IENA_MPRJ[92] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT37_A LA_DATA_OUT_CORE[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT380_A LA_IENA_MPRJ[93] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT381_A LA_IENA_MPRJ[94] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT382_A LA_IENA_MPRJ[95] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT383_A LA_IENA_MPRJ[96] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT384_A LA_IENA_MPRJ[97] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT385_A LA_IENA_MPRJ[98] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT386_A LA_IENA_MPRJ[99] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT387_A LA_IENA_MPRJ[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT388_A LA_OENB_MPRJ[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT389_A LA_OENB_MPRJ[100] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT38_A LA_DATA_OUT_CORE[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT390_A LA_OENB_MPRJ[101] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT391_A LA_OENB_MPRJ[102] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT392_A LA_OENB_MPRJ[103] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT393_A LA_OENB_MPRJ[104] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT394_A LA_OENB_MPRJ[105] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT395_A LA_OENB_MPRJ[106] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT396_A LA_OENB_MPRJ[107] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT397_A LA_OENB_MPRJ[108] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT398_A LA_OENB_MPRJ[109] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT399_A LA_OENB_MPRJ[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT39_A LA_DATA_OUT_CORE[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT3_A CARAVEL_RSTN VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT400_A LA_OENB_MPRJ[110] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT401_A LA_OENB_MPRJ[111] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT402_A LA_OENB_MPRJ[112] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT403_A LA_OENB_MPRJ[113] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT404_A LA_OENB_MPRJ[114] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT405_A LA_OENB_MPRJ[115] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT406_A LA_OENB_MPRJ[116] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT407_A LA_OENB_MPRJ[117] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT408_A LA_OENB_MPRJ[118] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT409_A LA_OENB_MPRJ[119] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT40_A LA_DATA_OUT_CORE[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT410_A LA_OENB_MPRJ[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT411_A LA_OENB_MPRJ[120] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT412_A LA_OENB_MPRJ[121] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT413_A LA_OENB_MPRJ[122] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT414_A LA_OENB_MPRJ[123] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT415_A LA_OENB_MPRJ[124] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT416_A LA_OENB_MPRJ[125] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT417_A LA_OENB_MPRJ[126] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT418_A LA_OENB_MPRJ[127] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT419_A LA_OENB_MPRJ[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT41_A LA_DATA_OUT_CORE[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT420_A LA_OENB_MPRJ[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT421_A LA_OENB_MPRJ[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT422_A LA_OENB_MPRJ[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT423_A LA_OENB_MPRJ[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT424_A LA_OENB_MPRJ[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT425_A LA_OENB_MPRJ[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT426_A LA_OENB_MPRJ[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT427_A LA_OENB_MPRJ[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT428_A LA_OENB_MPRJ[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT429_A LA_OENB_MPRJ[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT42_A LA_DATA_OUT_CORE[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT430_A LA_OENB_MPRJ[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT431_A LA_OENB_MPRJ[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT432_A LA_OENB_MPRJ[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT433_A LA_OENB_MPRJ[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT434_A LA_OENB_MPRJ[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT435_A LA_OENB_MPRJ[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT436_A LA_OENB_MPRJ[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT437_A LA_OENB_MPRJ[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT438_A LA_OENB_MPRJ[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT439_A LA_OENB_MPRJ[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT43_A LA_DATA_OUT_CORE[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT440_A LA_OENB_MPRJ[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT441_A LA_OENB_MPRJ[32] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT442_A LA_OENB_MPRJ[33] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT443_A LA_OENB_MPRJ[34] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT444_A LA_OENB_MPRJ[35] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT445_A LA_OENB_MPRJ[36] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT446_A LA_OENB_MPRJ[37] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT447_A LA_OENB_MPRJ[38] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT448_A LA_OENB_MPRJ[39] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT449_A LA_OENB_MPRJ[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT44_A LA_DATA_OUT_CORE[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT450_A LA_OENB_MPRJ[40] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT451_A LA_OENB_MPRJ[41] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT452_A LA_OENB_MPRJ[42] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT453_A LA_OENB_MPRJ[43] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT454_A LA_OENB_MPRJ[44] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT455_A LA_OENB_MPRJ[45] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT456_A LA_OENB_MPRJ[46] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT457_A LA_OENB_MPRJ[47] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT458_A LA_OENB_MPRJ[48] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT459_A LA_OENB_MPRJ[49] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT45_A LA_DATA_OUT_CORE[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT460_A LA_OENB_MPRJ[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT461_A LA_OENB_MPRJ[50] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT462_A LA_OENB_MPRJ[51] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT463_A LA_OENB_MPRJ[52] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT464_A LA_OENB_MPRJ[53] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT465_A LA_OENB_MPRJ[54] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT466_A LA_OENB_MPRJ[55] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT467_A LA_OENB_MPRJ[56] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT468_A LA_OENB_MPRJ[57] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT469_A LA_OENB_MPRJ[58] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT46_A LA_DATA_OUT_CORE[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT470_A LA_OENB_MPRJ[59] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT471_A LA_OENB_MPRJ[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT472_A LA_OENB_MPRJ[60] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT473_A LA_OENB_MPRJ[61] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT474_A LA_OENB_MPRJ[62] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT475_A LA_OENB_MPRJ[63] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT476_A LA_OENB_MPRJ[64] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT477_A LA_OENB_MPRJ[65] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT478_A LA_OENB_MPRJ[66] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT479_A LA_OENB_MPRJ[67] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT47_A LA_DATA_OUT_CORE[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT480_A LA_OENB_MPRJ[68] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT481_A LA_OENB_MPRJ[69] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT482_A LA_OENB_MPRJ[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT483_A LA_OENB_MPRJ[70] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT484_A LA_OENB_MPRJ[71] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT485_A LA_OENB_MPRJ[72] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT486_A LA_OENB_MPRJ[73] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT487_A LA_OENB_MPRJ[74] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT488_A LA_OENB_MPRJ[75] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT489_A LA_OENB_MPRJ[76] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT48_A LA_DATA_OUT_CORE[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT490_A LA_OENB_MPRJ[77] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT491_A LA_OENB_MPRJ[78] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT492_A LA_OENB_MPRJ[79] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT493_A LA_OENB_MPRJ[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT494_A LA_OENB_MPRJ[80] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT495_A LA_OENB_MPRJ[81] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT496_A LA_OENB_MPRJ[82] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT497_A LA_OENB_MPRJ[83] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT498_A LA_OENB_MPRJ[84] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT499_A LA_OENB_MPRJ[85] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT49_A LA_DATA_OUT_CORE[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT4_A LA_DATA_OUT_CORE[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT500_A LA_OENB_MPRJ[86] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT501_A LA_OENB_MPRJ[87] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT502_A LA_OENB_MPRJ[88] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT503_A LA_OENB_MPRJ[89] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT504_A LA_OENB_MPRJ[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT505_A LA_OENB_MPRJ[90] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT506_A LA_OENB_MPRJ[91] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT507_A LA_OENB_MPRJ[92] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT508_A LA_OENB_MPRJ[93] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT509_A LA_OENB_MPRJ[94] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT50_A LA_DATA_OUT_CORE[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT510_A LA_OENB_MPRJ[95] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT511_A LA_OENB_MPRJ[96] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT512_A LA_OENB_MPRJ[97] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT513_A LA_OENB_MPRJ[98] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT514_A LA_OENB_MPRJ[99] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT515_A LA_OENB_MPRJ[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT516_A MPRJ_ACK_I_USER VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT517_A MPRJ_ADR_O_CORE[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT518_A MPRJ_ADR_O_CORE[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT519_A MPRJ_ADR_O_CORE[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT51_A LA_DATA_OUT_CORE[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT520_A MPRJ_ADR_O_CORE[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT521_A MPRJ_ADR_O_CORE[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT522_A MPRJ_ADR_O_CORE[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT523_A MPRJ_ADR_O_CORE[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT524_A MPRJ_ADR_O_CORE[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT525_A MPRJ_ADR_O_CORE[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT526_A MPRJ_ADR_O_CORE[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT527_A MPRJ_ADR_O_CORE[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT528_A MPRJ_ADR_O_CORE[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT529_A MPRJ_ADR_O_CORE[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT52_A LA_DATA_OUT_CORE[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT530_A MPRJ_ADR_O_CORE[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT531_A MPRJ_ADR_O_CORE[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT532_A MPRJ_ADR_O_CORE[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT533_A MPRJ_ADR_O_CORE[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT534_A MPRJ_ADR_O_CORE[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT535_A MPRJ_ADR_O_CORE[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT536_A MPRJ_ADR_O_CORE[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT537_A MPRJ_ADR_O_CORE[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT538_A MPRJ_ADR_O_CORE[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT539_A MPRJ_ADR_O_CORE[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT53_A LA_DATA_OUT_CORE[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT540_A MPRJ_ADR_O_CORE[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT541_A MPRJ_ADR_O_CORE[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT542_A MPRJ_ADR_O_CORE[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT543_A MPRJ_ADR_O_CORE[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT544_A MPRJ_ADR_O_CORE[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT545_A MPRJ_ADR_O_CORE[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT546_A MPRJ_ADR_O_CORE[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT547_A MPRJ_ADR_O_CORE[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT548_A MPRJ_ADR_O_CORE[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT549_A MPRJ_CYC_O_CORE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT54_A LA_DATA_OUT_CORE[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT550_A MPRJ_DAT_I_USER[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT551_A MPRJ_DAT_I_USER[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT552_A MPRJ_DAT_I_USER[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT553_A MPRJ_DAT_I_USER[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT554_A MPRJ_DAT_I_USER[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT555_A MPRJ_DAT_I_USER[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT556_A MPRJ_DAT_I_USER[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT557_A MPRJ_DAT_I_USER[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT558_A MPRJ_DAT_I_USER[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT559_A MPRJ_DAT_I_USER[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT55_A LA_DATA_OUT_CORE[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT560_A MPRJ_DAT_I_USER[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT561_A MPRJ_DAT_I_USER[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT562_A MPRJ_DAT_I_USER[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT563_A MPRJ_DAT_I_USER[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT564_A MPRJ_DAT_I_USER[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT565_A MPRJ_DAT_I_USER[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT566_A MPRJ_DAT_I_USER[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT567_A MPRJ_DAT_I_USER[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT568_A MPRJ_DAT_I_USER[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT569_A MPRJ_DAT_I_USER[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT56_A LA_DATA_OUT_CORE[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT570_A MPRJ_DAT_I_USER[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT571_A MPRJ_DAT_I_USER[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT572_A MPRJ_DAT_I_USER[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT573_A MPRJ_DAT_I_USER[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT574_A MPRJ_DAT_I_USER[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT575_A MPRJ_DAT_I_USER[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT576_A MPRJ_DAT_I_USER[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT577_A MPRJ_DAT_I_USER[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT578_A MPRJ_DAT_I_USER[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT579_A MPRJ_DAT_I_USER[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT57_A LA_DATA_OUT_CORE[32] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT580_A MPRJ_DAT_I_USER[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT581_A MPRJ_DAT_I_USER[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT582_A MPRJ_DAT_O_CORE[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT583_A MPRJ_DAT_O_CORE[10] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT584_A MPRJ_DAT_O_CORE[11] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT585_A MPRJ_DAT_O_CORE[12] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT586_A MPRJ_DAT_O_CORE[13] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT587_A MPRJ_DAT_O_CORE[14] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT588_A MPRJ_DAT_O_CORE[15] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT589_A MPRJ_DAT_O_CORE[16] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT58_A LA_DATA_OUT_CORE[33] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT590_A MPRJ_DAT_O_CORE[17] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT591_A MPRJ_DAT_O_CORE[18] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT592_A MPRJ_DAT_O_CORE[19] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT593_A MPRJ_DAT_O_CORE[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT594_A MPRJ_DAT_O_CORE[20] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT595_A MPRJ_DAT_O_CORE[21] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT596_A MPRJ_DAT_O_CORE[22] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT597_A MPRJ_DAT_O_CORE[23] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT598_A MPRJ_DAT_O_CORE[24] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT599_A MPRJ_DAT_O_CORE[25] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT59_A LA_DATA_OUT_CORE[34] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT5_A LA_DATA_OUT_CORE[100] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT600_A MPRJ_DAT_O_CORE[26] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT601_A MPRJ_DAT_O_CORE[27] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT602_A MPRJ_DAT_O_CORE[28] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT603_A MPRJ_DAT_O_CORE[29] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT604_A MPRJ_DAT_O_CORE[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT605_A MPRJ_DAT_O_CORE[30] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT606_A MPRJ_DAT_O_CORE[31] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT607_A MPRJ_DAT_O_CORE[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT608_A MPRJ_DAT_O_CORE[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT609_A MPRJ_DAT_O_CORE[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT60_A LA_DATA_OUT_CORE[35] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT610_A MPRJ_DAT_O_CORE[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT611_A MPRJ_DAT_O_CORE[7] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT612_A MPRJ_DAT_O_CORE[8] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT613_A MPRJ_DAT_O_CORE[9] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT614_A MPRJ_IENA_WB VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT615_A MPRJ_SEL_O_CORE[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT616_A MPRJ_SEL_O_CORE[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT617_A MPRJ_SEL_O_CORE[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT618_A MPRJ_SEL_O_CORE[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT619_A MPRJ_STB_O_CORE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT61_A LA_DATA_OUT_CORE[36] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT620_A MPRJ_WE_O_CORE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT621_A USER_IRQ_CORE[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT622_A USER_IRQ_CORE[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT623_A USER_IRQ_CORE[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT624_A USER_IRQ_ENA[0] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT625_A USER_IRQ_ENA[1] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT626_A USER_IRQ_ENA[2] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT62_A LA_DATA_OUT_CORE[37] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT63_A LA_DATA_OUT_CORE[38] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT64_A LA_DATA_OUT_CORE[39] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT65_A LA_DATA_OUT_CORE[3] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT66_A LA_DATA_OUT_CORE[40] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT67_A LA_DATA_OUT_CORE[41] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT68_A LA_DATA_OUT_CORE[42] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT69_A LA_DATA_OUT_CORE[43] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT6_A LA_DATA_OUT_CORE[101] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT70_A LA_DATA_OUT_CORE[44] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT71_A LA_DATA_OUT_CORE[45] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT72_A LA_DATA_OUT_CORE[46] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT73_A LA_DATA_OUT_CORE[47] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT74_A LA_DATA_OUT_CORE[48] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT75_A LA_DATA_OUT_CORE[49] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT76_A LA_DATA_OUT_CORE[4] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT77_A LA_DATA_OUT_CORE[50] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT78_A LA_DATA_OUT_CORE[51] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT79_A LA_DATA_OUT_CORE[52] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT7_A LA_DATA_OUT_CORE[102] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT80_A LA_DATA_OUT_CORE[53] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT81_A LA_DATA_OUT_CORE[54] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT82_A LA_DATA_OUT_CORE[55] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT83_A LA_DATA_OUT_CORE[56] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT84_A LA_DATA_OUT_CORE[57] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT85_A LA_DATA_OUT_CORE[58] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT86_A LA_DATA_OUT_CORE[59] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT87_A LA_DATA_OUT_CORE[5] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT88_A LA_DATA_OUT_CORE[60] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT89_A LA_DATA_OUT_CORE[61] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT8_A LA_DATA_OUT_CORE[103] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT90_A LA_DATA_OUT_CORE[62] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT91_A LA_DATA_OUT_CORE[63] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT92_A LA_DATA_OUT_CORE[64] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT93_A LA_DATA_OUT_CORE[65] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT94_A LA_DATA_OUT_CORE[66] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT95_A LA_DATA_OUT_CORE[67] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT96_A LA_DATA_OUT_CORE[68] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT97_A LA_DATA_OUT_CORE[69] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT98_A LA_DATA_OUT_CORE[6] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT99_A LA_DATA_OUT_CORE[70] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_INPUT9_A LA_DATA_OUT_CORE[104] VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[0]_A _073_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[0]_TE \LA_DATA_OUT_ENABLE[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[100]_A _074_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[100]_TE \LA_DATA_OUT_ENABLE[100]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[101]_A _075_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[101]_TE \LA_DATA_OUT_ENABLE[101]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[102]_A _076_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[102]_TE \LA_DATA_OUT_ENABLE[102]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[103]_A _077_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[103]_TE \LA_DATA_OUT_ENABLE[103]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[104]_A _078_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[104]_TE \LA_DATA_OUT_ENABLE[104]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[105]_A _079_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[105]_TE \LA_DATA_OUT_ENABLE[105]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[106]_A _080_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[106]_TE \LA_DATA_OUT_ENABLE[106]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[107]_A _081_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[107]_TE \LA_DATA_OUT_ENABLE[107]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[108]_A _082_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[108]_TE \LA_DATA_OUT_ENABLE[108]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[109]_A _083_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[109]_TE \LA_DATA_OUT_ENABLE[109]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[10]_A _084_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[10]_TE \LA_DATA_OUT_ENABLE[10]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[110]_A _085_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[110]_TE \LA_DATA_OUT_ENABLE[110]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[111]_A _086_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[111]_TE \LA_DATA_OUT_ENABLE[111]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[112]_A _087_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[112]_TE \LA_DATA_OUT_ENABLE[112]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[113]_A _088_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[113]_TE \LA_DATA_OUT_ENABLE[113]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[114]_A _089_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[114]_TE \LA_DATA_OUT_ENABLE[114]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[115]_A _090_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[115]_TE \LA_DATA_OUT_ENABLE[115]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[116]_A _091_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[116]_TE \LA_DATA_OUT_ENABLE[116]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[117]_A _092_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[117]_TE \LA_DATA_OUT_ENABLE[117]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[118]_A _093_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[118]_TE \LA_DATA_OUT_ENABLE[118]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[119]_A _094_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[119]_TE \LA_DATA_OUT_ENABLE[119]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[11]_A _095_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[11]_TE \LA_DATA_OUT_ENABLE[11]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[120]_A _096_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[120]_TE \LA_DATA_OUT_ENABLE[120]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[121]_A _097_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[121]_TE \LA_DATA_OUT_ENABLE[121]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[122]_A _098_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[122]_TE \LA_DATA_OUT_ENABLE[122]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[123]_A _099_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[123]_TE \LA_DATA_OUT_ENABLE[123]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[124]_A _100_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[124]_TE \LA_DATA_OUT_ENABLE[124]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[125]_A _101_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[125]_TE \LA_DATA_OUT_ENABLE[125]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[126]_A _102_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[126]_TE \LA_DATA_OUT_ENABLE[126]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[127]_A _103_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[127]_TE \LA_DATA_OUT_ENABLE[127]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[12]_A _104_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[12]_TE \LA_DATA_OUT_ENABLE[12]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[13]_A _105_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[13]_TE \LA_DATA_OUT_ENABLE[13]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[14]_A _106_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[14]_TE \LA_DATA_OUT_ENABLE[14]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[15]_A _107_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[15]_TE \LA_DATA_OUT_ENABLE[15]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[16]_A _108_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[16]_TE \LA_DATA_OUT_ENABLE[16]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[17]_A _109_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[17]_TE \LA_DATA_OUT_ENABLE[17]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[18]_A _110_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[18]_TE \LA_DATA_OUT_ENABLE[18]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[19]_A _111_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[19]_TE \LA_DATA_OUT_ENABLE[19]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[1]_A _112_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[1]_TE \LA_DATA_OUT_ENABLE[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[20]_A _113_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[20]_TE \LA_DATA_OUT_ENABLE[20]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[21]_A _114_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[21]_TE \LA_DATA_OUT_ENABLE[21]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[22]_A _115_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[22]_TE \LA_DATA_OUT_ENABLE[22]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[23]_A _116_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[23]_TE \LA_DATA_OUT_ENABLE[23]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[24]_A _117_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[24]_TE \LA_DATA_OUT_ENABLE[24]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[25]_A _118_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[25]_TE \LA_DATA_OUT_ENABLE[25]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[26]_A _119_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[26]_TE \LA_DATA_OUT_ENABLE[26]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[27]_A _120_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[27]_TE \LA_DATA_OUT_ENABLE[27]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[28]_A _121_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[28]_TE \LA_DATA_OUT_ENABLE[28]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[29]_A _122_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[29]_TE \LA_DATA_OUT_ENABLE[29]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[2]_A _123_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[2]_TE \LA_DATA_OUT_ENABLE[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[30]_A _124_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[30]_TE \LA_DATA_OUT_ENABLE[30]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[31]_A _125_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[31]_TE \LA_DATA_OUT_ENABLE[31]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[32]_A _126_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[32]_TE \LA_DATA_OUT_ENABLE[32]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[33]_A _127_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[33]_TE \LA_DATA_OUT_ENABLE[33]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[34]_A _128_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[34]_TE \LA_DATA_OUT_ENABLE[34]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[35]_A _129_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[35]_TE \LA_DATA_OUT_ENABLE[35]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[36]_A _130_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[36]_TE \LA_DATA_OUT_ENABLE[36]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[37]_A _131_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[37]_TE \LA_DATA_OUT_ENABLE[37]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[38]_A _132_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[38]_TE \LA_DATA_OUT_ENABLE[38]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[39]_A _133_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[39]_TE \LA_DATA_OUT_ENABLE[39]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[3]_A _134_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[3]_TE \LA_DATA_OUT_ENABLE[3]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[40]_A _135_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[40]_TE \LA_DATA_OUT_ENABLE[40]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[41]_A _136_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[41]_TE \LA_DATA_OUT_ENABLE[41]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[42]_A _137_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[42]_TE \LA_DATA_OUT_ENABLE[42]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[43]_A _138_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[43]_TE \LA_DATA_OUT_ENABLE[43]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[44]_A _139_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[44]_TE \LA_DATA_OUT_ENABLE[44]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[45]_A _140_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[45]_TE \LA_DATA_OUT_ENABLE[45]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[46]_A _141_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[46]_TE \LA_DATA_OUT_ENABLE[46]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[47]_A _142_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[47]_TE \LA_DATA_OUT_ENABLE[47]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[48]_A _143_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[48]_TE \LA_DATA_OUT_ENABLE[48]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[49]_A _144_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[49]_TE \LA_DATA_OUT_ENABLE[49]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[4]_A _145_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[4]_TE \LA_DATA_OUT_ENABLE[4]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[50]_A _146_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[50]_TE \LA_DATA_OUT_ENABLE[50]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[51]_A _147_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[51]_TE \LA_DATA_OUT_ENABLE[51]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[52]_A _148_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[52]_TE \LA_DATA_OUT_ENABLE[52]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[53]_A _149_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[53]_TE \LA_DATA_OUT_ENABLE[53]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[54]_A _150_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[54]_TE \LA_DATA_OUT_ENABLE[54]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[55]_A _151_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[55]_TE \LA_DATA_OUT_ENABLE[55]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[56]_A _152_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[56]_TE \LA_DATA_OUT_ENABLE[56]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[57]_A _153_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[57]_TE \LA_DATA_OUT_ENABLE[57]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[58]_A _154_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[58]_TE \LA_DATA_OUT_ENABLE[58]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[59]_A _155_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[59]_TE \LA_DATA_OUT_ENABLE[59]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[5]_A _156_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[5]_TE \LA_DATA_OUT_ENABLE[5]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[60]_A _157_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[60]_TE \LA_DATA_OUT_ENABLE[60]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[61]_A _158_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[61]_TE \LA_DATA_OUT_ENABLE[61]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[62]_A _159_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[62]_TE \LA_DATA_OUT_ENABLE[62]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[63]_A _160_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[63]_TE \LA_DATA_OUT_ENABLE[63]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[64]_A _161_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[64]_TE \LA_DATA_OUT_ENABLE[64]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[65]_A _162_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[65]_TE \LA_DATA_OUT_ENABLE[65]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[66]_A _163_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[66]_TE \LA_DATA_OUT_ENABLE[66]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[67]_A _164_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[67]_TE \LA_DATA_OUT_ENABLE[67]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[68]_A _165_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[68]_TE \LA_DATA_OUT_ENABLE[68]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[69]_A _166_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[69]_TE \LA_DATA_OUT_ENABLE[69]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[6]_A _167_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[6]_TE \LA_DATA_OUT_ENABLE[6]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[70]_A _168_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[70]_TE \LA_DATA_OUT_ENABLE[70]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[71]_A _169_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[71]_TE \LA_DATA_OUT_ENABLE[71]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[72]_A _170_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[72]_TE \LA_DATA_OUT_ENABLE[72]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[73]_A _171_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[73]_TE \LA_DATA_OUT_ENABLE[73]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[74]_A _172_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[74]_TE \LA_DATA_OUT_ENABLE[74]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[75]_A _173_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[75]_TE \LA_DATA_OUT_ENABLE[75]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[76]_A _174_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[76]_TE \LA_DATA_OUT_ENABLE[76]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[77]_A _175_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[77]_TE \LA_DATA_OUT_ENABLE[77]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[78]_A _176_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[78]_TE \LA_DATA_OUT_ENABLE[78]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[79]_A _177_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[79]_TE \LA_DATA_OUT_ENABLE[79]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[7]_A _178_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[7]_TE \LA_DATA_OUT_ENABLE[7]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[80]_A _179_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[80]_TE \LA_DATA_OUT_ENABLE[80]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[81]_A _180_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[81]_TE \LA_DATA_OUT_ENABLE[81]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[82]_A _181_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[82]_TE \LA_DATA_OUT_ENABLE[82]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[83]_A _182_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[83]_TE \LA_DATA_OUT_ENABLE[83]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[84]_A _183_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[84]_TE \LA_DATA_OUT_ENABLE[84]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[85]_A _184_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[85]_TE \LA_DATA_OUT_ENABLE[85]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[86]_A _185_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[86]_TE \LA_DATA_OUT_ENABLE[86]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[87]_A _186_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[87]_TE \LA_DATA_OUT_ENABLE[87]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[88]_A _187_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[88]_TE \LA_DATA_OUT_ENABLE[88]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[89]_A _188_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[89]_TE \LA_DATA_OUT_ENABLE[89]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[8]_A _189_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[8]_TE \LA_DATA_OUT_ENABLE[8]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[90]_A _190_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[90]_TE \LA_DATA_OUT_ENABLE[90]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[91]_A _191_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[91]_TE \LA_DATA_OUT_ENABLE[91]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[92]_A _192_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[92]_TE \LA_DATA_OUT_ENABLE[92]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[93]_A _193_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[93]_TE \LA_DATA_OUT_ENABLE[93]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[94]_A _194_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[94]_TE \LA_DATA_OUT_ENABLE[94]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[95]_A _195_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[95]_TE \LA_DATA_OUT_ENABLE[95]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[96]_A _196_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[96]_TE \LA_DATA_OUT_ENABLE[96]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[97]_A _197_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[97]_TE \LA_DATA_OUT_ENABLE[97]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[98]_A _198_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[98]_TE \LA_DATA_OUT_ENABLE[98]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[99]_A _199_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[99]_TE \LA_DATA_OUT_ENABLE[99]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[9]_A _200_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF[9]_TE \LA_DATA_OUT_ENABLE[9]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[0]_A_N NET388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[0]_B \MPRJ_LOGIC1[74]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[100]_A_N NET389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[100]_B \MPRJ_LOGIC1[174]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[101]_A_N NET390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[101]_B \MPRJ_LOGIC1[175]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[102]_A_N NET391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[102]_B \MPRJ_LOGIC1[176]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[103]_A_N NET392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[103]_B \MPRJ_LOGIC1[177]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[104]_A_N NET393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[104]_B \MPRJ_LOGIC1[178]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[105]_A_N NET394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[105]_B \MPRJ_LOGIC1[179]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[106]_A_N NET395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[106]_B \MPRJ_LOGIC1[180]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[107]_A_N NET396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[107]_B \MPRJ_LOGIC1[181]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[108]_A_N NET397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[108]_B \MPRJ_LOGIC1[182]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[109]_A_N NET398 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[109]_B \MPRJ_LOGIC1[183]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[10]_A_N NET399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[10]_B \MPRJ_LOGIC1[84]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[110]_A_N NET400 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[110]_B \MPRJ_LOGIC1[184]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[111]_A_N NET401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[111]_B \MPRJ_LOGIC1[185]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[112]_A_N NET402 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[112]_B \MPRJ_LOGIC1[186]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[113]_A_N NET403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[113]_B \MPRJ_LOGIC1[187]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[114]_A_N NET404 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[114]_B \MPRJ_LOGIC1[188]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[115]_A_N NET405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[115]_B \MPRJ_LOGIC1[189]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[116]_A_N NET406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[116]_B \MPRJ_LOGIC1[190]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[117]_A_N NET407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[117]_B \MPRJ_LOGIC1[191]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[118]_A_N NET408 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[118]_B \MPRJ_LOGIC1[192]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[119]_A_N NET409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[119]_B \MPRJ_LOGIC1[193]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[11]_A_N NET410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[11]_B \MPRJ_LOGIC1[85]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[120]_A_N NET411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[120]_B \MPRJ_LOGIC1[194]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[121]_A_N NET412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[121]_B \MPRJ_LOGIC1[195]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[122]_A_N NET413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[122]_B \MPRJ_LOGIC1[196]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[123]_A_N NET414 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[123]_B \MPRJ_LOGIC1[197]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[124]_A_N NET415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[124]_B \MPRJ_LOGIC1[198]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[125]_A_N NET416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[125]_B \MPRJ_LOGIC1[199]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[126]_A_N NET417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[126]_B \MPRJ_LOGIC1[200]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[127]_A_N NET418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[127]_B \MPRJ_LOGIC1[201]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[12]_A_N NET419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[12]_B \MPRJ_LOGIC1[86]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[13]_A_N NET420 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[13]_B \MPRJ_LOGIC1[87]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[14]_A_N NET421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[14]_B \MPRJ_LOGIC1[88]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[15]_A_N NET422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[15]_B \MPRJ_LOGIC1[89]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[16]_A_N NET423 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[16]_B \MPRJ_LOGIC1[90]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[17]_A_N NET424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[17]_B \MPRJ_LOGIC1[91]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[18]_A_N NET425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[18]_B \MPRJ_LOGIC1[92]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[19]_A_N NET426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[19]_B \MPRJ_LOGIC1[93]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[1]_A_N NET427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[1]_B \MPRJ_LOGIC1[75]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[20]_A_N NET428 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[20]_B \MPRJ_LOGIC1[94]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[21]_A_N NET429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[21]_B \MPRJ_LOGIC1[95]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[22]_A_N NET430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[22]_B \MPRJ_LOGIC1[96]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[23]_A_N NET431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[23]_B \MPRJ_LOGIC1[97]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[24]_A_N NET432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[24]_B \MPRJ_LOGIC1[98]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[25]_A_N NET433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[25]_B \MPRJ_LOGIC1[99]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[26]_A_N NET434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[26]_B \MPRJ_LOGIC1[100]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[27]_A_N NET435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[27]_B \MPRJ_LOGIC1[101]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[28]_A_N NET436 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[28]_B \MPRJ_LOGIC1[102]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[29]_A_N NET437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[29]_B \MPRJ_LOGIC1[103]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[2]_A_N NET438 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[2]_B \MPRJ_LOGIC1[76]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[30]_A_N NET439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[30]_B \MPRJ_LOGIC1[104]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[31]_A_N NET440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[31]_B \MPRJ_LOGIC1[105]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[32]_A_N NET441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[32]_B \MPRJ_LOGIC1[106]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[33]_A_N NET442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[33]_B \MPRJ_LOGIC1[107]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[34]_A_N NET443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[34]_B \MPRJ_LOGIC1[108]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[35]_A_N NET444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[35]_B \MPRJ_LOGIC1[109]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[36]_A_N NET445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[36]_B \MPRJ_LOGIC1[110]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[37]_A_N NET446 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[37]_B \MPRJ_LOGIC1[111]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[38]_A_N NET447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[38]_B \MPRJ_LOGIC1[112]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[39]_A_N NET448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[39]_B \MPRJ_LOGIC1[113]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[3]_A_N NET449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[3]_B \MPRJ_LOGIC1[77]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[40]_A_N NET450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[40]_B \MPRJ_LOGIC1[114]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[41]_A_N NET451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[41]_B \MPRJ_LOGIC1[115]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[42]_A_N NET452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[42]_B \MPRJ_LOGIC1[116]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[43]_A_N NET453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[43]_B \MPRJ_LOGIC1[117]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[44]_A_N NET454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[44]_B \MPRJ_LOGIC1[118]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[45]_A_N NET455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[45]_B \MPRJ_LOGIC1[119]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[46]_A_N NET456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[46]_B \MPRJ_LOGIC1[120]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[47]_A_N NET457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[47]_B \MPRJ_LOGIC1[121]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[48]_A_N NET458 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[48]_B \MPRJ_LOGIC1[122]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[49]_A_N NET459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[49]_B \MPRJ_LOGIC1[123]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[4]_A_N NET460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[4]_B \MPRJ_LOGIC1[78]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[50]_A_N NET461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[50]_B \MPRJ_LOGIC1[124]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[51]_A_N NET462 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[51]_B \MPRJ_LOGIC1[125]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[52]_A_N NET463 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[52]_B \MPRJ_LOGIC1[126]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[53]_A_N NET464 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[53]_B \MPRJ_LOGIC1[127]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[54]_A_N NET465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[54]_B \MPRJ_LOGIC1[128]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[55]_A_N NET466 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[55]_B \MPRJ_LOGIC1[129]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[56]_A_N NET467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[56]_B \MPRJ_LOGIC1[130]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[57]_A_N NET468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[57]_B \MPRJ_LOGIC1[131]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[58]_A_N NET469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[58]_B \MPRJ_LOGIC1[132]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[59]_A_N NET470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[59]_B \MPRJ_LOGIC1[133]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[5]_A_N NET471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[5]_B \MPRJ_LOGIC1[79]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[60]_A_N NET472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[60]_B \MPRJ_LOGIC1[134]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[61]_A_N NET473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[61]_B \MPRJ_LOGIC1[135]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[62]_A_N NET474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[62]_B \MPRJ_LOGIC1[136]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[63]_A_N NET475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[63]_B \MPRJ_LOGIC1[137]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[64]_A_N NET476 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[64]_B \MPRJ_LOGIC1[138]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[65]_A_N NET477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[65]_B \MPRJ_LOGIC1[139]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[66]_A_N NET478 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[66]_B \MPRJ_LOGIC1[140]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[67]_A_N NET479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[67]_B \MPRJ_LOGIC1[141]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[68]_A_N NET480 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[68]_B \MPRJ_LOGIC1[142]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[69]_A_N NET481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[69]_B \MPRJ_LOGIC1[143]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[6]_A_N NET482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[6]_B \MPRJ_LOGIC1[80]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[70]_A_N NET483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[70]_B \MPRJ_LOGIC1[144]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[71]_A_N NET484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[71]_B \MPRJ_LOGIC1[145]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[72]_A_N NET485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[72]_B \MPRJ_LOGIC1[146]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[73]_A_N NET486 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[73]_B \MPRJ_LOGIC1[147]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[74]_A_N NET487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[74]_B \MPRJ_LOGIC1[148]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[75]_A_N NET488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[75]_B \MPRJ_LOGIC1[149]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[76]_A_N NET489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[76]_B \MPRJ_LOGIC1[150]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[77]_A_N NET490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[77]_B \MPRJ_LOGIC1[151]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[78]_A_N NET491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[78]_B \MPRJ_LOGIC1[152]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[79]_A_N NET492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[79]_B \MPRJ_LOGIC1[153]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[7]_A_N NET493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[7]_B \MPRJ_LOGIC1[81]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[80]_A_N NET494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[80]_B \MPRJ_LOGIC1[154]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[81]_A_N NET495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[81]_B \MPRJ_LOGIC1[155]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[82]_A_N NET496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[82]_B \MPRJ_LOGIC1[156]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[83]_A_N NET497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[83]_B \MPRJ_LOGIC1[157]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[84]_A_N NET498 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[84]_B \MPRJ_LOGIC1[158]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[85]_A_N NET499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[85]_B \MPRJ_LOGIC1[159]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[86]_A_N NET500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[86]_B \MPRJ_LOGIC1[160]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[87]_A_N NET501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[87]_B \MPRJ_LOGIC1[161]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[88]_A_N NET502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[88]_B \MPRJ_LOGIC1[162]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[89]_A_N NET503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[89]_B \MPRJ_LOGIC1[163]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[8]_A_N NET504 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[8]_B \MPRJ_LOGIC1[82]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[90]_A_N NET505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[90]_B \MPRJ_LOGIC1[164]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[91]_A_N NET506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[91]_B \MPRJ_LOGIC1[165]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[92]_A_N NET507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[92]_B \MPRJ_LOGIC1[166]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[93]_A_N NET508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[93]_B \MPRJ_LOGIC1[167]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[94]_A_N NET509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[94]_B \MPRJ_LOGIC1[168]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[95]_A_N NET510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[95]_B \MPRJ_LOGIC1[169]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[96]_A_N NET511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[96]_B \MPRJ_LOGIC1[170]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[97]_A_N NET512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[97]_B \MPRJ_LOGIC1[171]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[98]_A_N NET513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[98]_B \MPRJ_LOGIC1[172]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[99]_A_N NET514 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[99]_B \MPRJ_LOGIC1[173]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[9]_A_N NET515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_LA_BUF_ENABLE[9]_B \MPRJ_LOGIC1[83]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ2_PWRGOOD_A MPRJ2_LOGIC1 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ2_VDD_PWRGOOD_A MPRJ2_VDD_LOGIC1 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[0]_A _009_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[0]_TE \MPRJ_LOGIC1[10]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[10]_A _010_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[10]_TE \MPRJ_LOGIC1[20]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[11]_A _011_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[11]_TE \MPRJ_LOGIC1[21]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[12]_A _012_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[12]_TE \MPRJ_LOGIC1[22]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[13]_A _013_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[13]_TE \MPRJ_LOGIC1[23]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[14]_A _014_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[14]_TE \MPRJ_LOGIC1[24]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[15]_A _015_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[15]_TE \MPRJ_LOGIC1[25]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[16]_A _016_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[16]_TE \MPRJ_LOGIC1[26]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[17]_A _017_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[17]_TE \MPRJ_LOGIC1[27]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[18]_A _018_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[18]_TE \MPRJ_LOGIC1[28]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[19]_A _019_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[19]_TE \MPRJ_LOGIC1[29]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[1]_A _020_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[1]_TE \MPRJ_LOGIC1[11]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[20]_A _021_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[20]_TE \MPRJ_LOGIC1[30]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[21]_A _022_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[21]_TE \MPRJ_LOGIC1[31]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[22]_A _023_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[22]_TE \MPRJ_LOGIC1[32]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[23]_A _024_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[23]_TE \MPRJ_LOGIC1[33]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[24]_A _025_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[24]_TE \MPRJ_LOGIC1[34]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[25]_A _026_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[25]_TE \MPRJ_LOGIC1[35]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[26]_A _027_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[26]_TE \MPRJ_LOGIC1[36]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[27]_A _028_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[27]_TE \MPRJ_LOGIC1[37]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[28]_A _029_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[28]_TE \MPRJ_LOGIC1[38]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[29]_A _030_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[29]_TE \MPRJ_LOGIC1[39]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[2]_A _031_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[2]_TE \MPRJ_LOGIC1[12]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[30]_A _032_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[30]_TE \MPRJ_LOGIC1[40]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[31]_A _033_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[31]_TE \MPRJ_LOGIC1[41]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[3]_A _034_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[3]_TE \MPRJ_LOGIC1[13]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[4]_A _035_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[4]_TE \MPRJ_LOGIC1[14]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[5]_A _036_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[5]_TE \MPRJ_LOGIC1[15]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[6]_A _037_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[6]_TE \MPRJ_LOGIC1[16]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[7]_A _038_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[7]_TE \MPRJ_LOGIC1[17]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[8]_A _039_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[8]_TE \MPRJ_LOGIC1[18]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[9]_A _040_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_ADR_BUF[9]_TE \MPRJ_LOGIC1[19]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CLK2_BUF_A _001_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CLK2_BUF_TE \MPRJ_LOGIC1[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CLK_BUF_A _000_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CLK_BUF_TE \MPRJ_LOGIC1[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CYC_BUF_A _002_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_CYC_BUF_TE \MPRJ_LOGIC1[3]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[0]_A _041_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[0]_TE \MPRJ_LOGIC1[42]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[10]_A _042_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[10]_TE \MPRJ_LOGIC1[52]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[11]_A _043_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[11]_TE \MPRJ_LOGIC1[53]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[12]_A _044_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[12]_TE \MPRJ_LOGIC1[54]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[13]_A _045_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[13]_TE \MPRJ_LOGIC1[55]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[14]_A _046_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[14]_TE \MPRJ_LOGIC1[56]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[15]_A _047_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[15]_TE \MPRJ_LOGIC1[57]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[16]_A _048_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[16]_TE \MPRJ_LOGIC1[58]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[17]_A _049_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[17]_TE \MPRJ_LOGIC1[59]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[18]_A _050_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[18]_TE \MPRJ_LOGIC1[60]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[19]_A _051_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[19]_TE \MPRJ_LOGIC1[61]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[1]_A _052_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[1]_TE \MPRJ_LOGIC1[43]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[20]_A _053_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[20]_TE \MPRJ_LOGIC1[62]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[21]_A _054_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[21]_TE \MPRJ_LOGIC1[63]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[22]_A _055_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[22]_TE \MPRJ_LOGIC1[64]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[23]_A _056_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[23]_TE \MPRJ_LOGIC1[65]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[24]_A _057_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[24]_TE \MPRJ_LOGIC1[66]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[25]_A _058_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[25]_TE \MPRJ_LOGIC1[67]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[26]_A _059_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[26]_TE \MPRJ_LOGIC1[68]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[27]_A _060_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[27]_TE \MPRJ_LOGIC1[69]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[28]_A _061_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[28]_TE \MPRJ_LOGIC1[70]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[29]_A _062_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[29]_TE \MPRJ_LOGIC1[71]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[2]_A _063_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[2]_TE \MPRJ_LOGIC1[44]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[30]_A _064_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[30]_TE \MPRJ_LOGIC1[72]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[31]_A _065_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[31]_TE \MPRJ_LOGIC1[73]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[3]_A _066_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[3]_TE \MPRJ_LOGIC1[45]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[4]_A _067_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[4]_TE \MPRJ_LOGIC1[46]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[5]_A _068_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[5]_TE \MPRJ_LOGIC1[47]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[6]_A _069_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[6]_TE \MPRJ_LOGIC1[48]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[7]_A _070_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[7]_TE \MPRJ_LOGIC1[49]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[8]_A _071_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[8]_TE \MPRJ_LOGIC1[50]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[9]_A _072_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_DAT_BUF[9]_TE \MPRJ_LOGIC1[51]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_PWRGOOD_A \MPRJ_LOGIC1[461]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_RSTN_BUF_A NET3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_RSTN_BUF_TE \MPRJ_LOGIC1[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[0]_A _005_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[0]_TE \MPRJ_LOGIC1[6]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[1]_A _006_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[1]_TE \MPRJ_LOGIC1[7]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[2]_A _007_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[2]_TE \MPRJ_LOGIC1[8]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[3]_A _008_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_MPRJ_SEL_BUF[3]_TE \MPRJ_LOGIC1[9]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_STB_BUF_A _003_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_STB_BUF_TE \MPRJ_LOGIC1[4]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_VDD_PWRGOOD_A MPRJ_VDD_LOGIC1 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_WE_BUF_A _004_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_MPRJ_WE_BUF_TE \MPRJ_LOGIC1[5]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1000_A NET1000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1001_A NET1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1002_A NET1002 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1003_A NET1003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1004_A NET1004 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1005_A NET1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1006_A NET1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1007_A NET1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1008_A NET1008 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1009_A NET1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1010_A NET1010 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1011_A NET1011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1012_A NET1012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1013_A NET1013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1014_A NET1014 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1015_A NET1015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1016_A NET1016 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1017_A NET1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1018_A NET1018 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1019_A NET1019 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1020_A NET1020 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1021_A NET1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1022_A NET1022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1023_A NET1023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1024_A NET1024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1025_A NET1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1026_A NET1026 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1027_A NET1027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1028_A NET1028 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1029_A NET1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1030_A NET1030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1031_A NET1031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1032_A NET1032 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1033_A NET1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1034_A NET1034 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1035_A NET1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1036_A NET1036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1037_A NET1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1038_A NET1038 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1039_A NET1039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1040_A NET1040 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1041_A NET1041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1042_A NET1042 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1043_A NET1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1044_A NET1044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1045_A NET1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1046_A NET1046 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1047_A NET1047 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1048_A NET1048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1049_A NET1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1050_A NET1050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1051_A NET1051 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1052_A NET1052 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1053_A NET1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1054_A NET1054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1055_A NET1055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1056_A NET1056 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1057_A NET1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1058_A NET1058 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1059_A NET1059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1060_A NET1060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1061_A NET1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1062_A NET1062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1063_A NET1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1064_A NET1064 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1065_A NET1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1066_A NET1066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1067_A NET1067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1068_A NET1068 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1069_A NET1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1070_A NET1070 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1071_A NET1071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1072_A NET1072 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1073_A NET1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1074_A NET1074 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1075_A NET1075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1076_A NET1076 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1077_A NET1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1078_A NET1078 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1079_A NET1079 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1080_A NET1080 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1081_A NET1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1082_A NET1082 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1083_A NET1083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1084_A NET1084 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1085_A NET1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1086_A NET1086 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1087_A NET1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1088_A NET1088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1089_A NET1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1090_A NET1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1091_A NET1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1092_A NET1092 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1093_A NET1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1094_A NET1094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1095_A NET1095 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1096_A NET1096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1097_A NET1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1098_A NET1098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1099_A NET1099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1100_A NET1100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1101_A NET1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1102_A NET1102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1103_A NET1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1104_A NET1104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1105_A NET1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1106_A NET1106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1107_A NET1107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1108_A NET1108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1109_A NET1109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1110_A NET1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1111_A NET1111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1112_A NET1112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1113_A NET1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1114_A NET1114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1115_A NET1115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1116_A NET1116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1117_A NET1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1118_A NET1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1119_A NET1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1120_A NET1120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1121_A NET1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1122_A NET1122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1123_A NET1123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT1124_A NET1124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT627_A NET627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT628_A NET628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT629_A NET629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT630_A NET630 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT631_A NET631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT632_A NET632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT633_A NET633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT634_A NET634 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT635_A NET635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT636_A NET636 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT637_A NET637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT638_A NET638 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT639_A NET639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT640_A NET640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT641_A NET641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT642_A NET642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT643_A NET643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT644_A NET644 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT645_A NET645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT646_A NET646 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT647_A NET647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT648_A NET648 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT649_A NET649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT650_A NET650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT651_A NET651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT652_A NET652 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT653_A NET653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT654_A NET654 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT655_A NET655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT656_A NET656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT657_A NET657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT658_A NET658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT659_A NET659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT660_A NET660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT661_A NET661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT662_A NET662 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT663_A NET663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT664_A NET664 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT665_A NET665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT666_A NET666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT667_A NET667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT668_A NET668 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT669_A NET669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT670_A NET670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT671_A NET671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT672_A NET672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT673_A NET673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT674_A NET674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT675_A NET675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT676_A NET676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT677_A NET677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT678_A NET678 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT679_A NET679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT680_A NET680 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT681_A NET681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT682_A NET682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT683_A NET683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT684_A NET684 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT685_A NET685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT686_A NET686 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT687_A NET687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT688_A NET688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT689_A NET689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT690_A NET690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT691_A NET691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT692_A NET692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT693_A NET693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT694_A NET694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT695_A NET695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT696_A NET696 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT697_A NET697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT698_A NET698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT699_A NET699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT700_A NET700 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT701_A NET701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT702_A NET702 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT703_A NET703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT704_A NET704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT705_A NET705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT706_A NET706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT707_A NET707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT708_A NET708 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT709_A NET709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT710_A NET710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT711_A NET711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT712_A NET712 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT713_A NET713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT714_A NET714 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT715_A NET715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT716_A NET716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT717_A NET717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT718_A NET718 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT719_A NET719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT720_A NET720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT721_A NET721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT722_A NET722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT723_A NET723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT724_A NET724 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT725_A NET725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT726_A NET726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT727_A NET727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT728_A NET728 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT729_A NET729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT730_A NET730 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT731_A NET731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT732_A NET732 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT733_A NET733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT734_A NET734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT735_A NET735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT736_A NET736 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT737_A NET737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT738_A NET738 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT739_A NET739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT740_A NET740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT741_A NET741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT742_A NET742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT743_A NET743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT744_A NET744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT745_A NET745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT746_A NET746 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT747_A NET747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT748_A NET748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT749_A NET749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT750_A NET750 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT751_A NET751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT752_A NET752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT753_A NET753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT754_A NET754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT755_A NET755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT756_A NET756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT757_A NET757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT758_A NET758 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT759_A NET759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT760_A NET760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT761_A NET761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT762_A NET762 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT763_A NET763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT764_A NET764 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT765_A NET765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT766_A NET766 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT767_A NET767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT768_A NET768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT769_A NET769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT770_A NET770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT771_A NET771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT772_A NET772 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT773_A NET773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT774_A NET774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT775_A NET775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT776_A NET776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT777_A NET777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT778_A NET778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT779_A NET779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT780_A NET780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT781_A NET781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT782_A NET782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT783_A NET783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT784_A NET784 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT785_A NET785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT786_A NET786 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT787_A NET787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT788_A NET788 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT789_A NET789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT790_A NET790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT791_A NET791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT792_A NET792 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT793_A NET793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT794_A NET794 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT795_A NET795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT796_A NET796 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT797_A NET797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT798_A NET798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT799_A NET799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT800_A NET800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT801_A NET801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT802_A NET802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT803_A NET803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT804_A NET804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT805_A NET805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT806_A NET806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT807_A NET807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT808_A NET808 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT809_A NET809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT810_A NET810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT811_A NET811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT812_A NET812 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT813_A NET813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT814_A NET814 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT815_A NET815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT816_A NET816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT817_A NET817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT818_A NET818 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT819_A NET819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT820_A NET820 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT821_A NET821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT822_A NET822 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT823_A NET823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT824_A NET824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT825_A NET825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT826_A NET826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT827_A NET827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT828_A NET828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT829_A NET829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT830_A NET830 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT831_A NET831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT832_A NET832 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT833_A NET833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT834_A NET834 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT835_A NET835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT836_A NET836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT837_A NET837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT838_A NET838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT839_A NET839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT840_A NET840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT841_A NET841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT842_A NET842 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT843_A NET843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT844_A NET844 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT845_A NET845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT846_A NET846 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT847_A NET847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT848_A NET848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT849_A NET849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT850_A NET850 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT851_A NET851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT852_A NET852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT853_A NET853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT854_A NET854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT855_A NET855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT856_A NET856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT857_A NET857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT858_A NET858 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT859_A NET859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT860_A NET860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT861_A NET861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT862_A NET862 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT863_A NET863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT864_A NET864 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT865_A NET865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT866_A NET866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT867_A NET867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT868_A NET868 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT869_A NET869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT870_A NET870 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT871_A NET871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT872_A NET872 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT873_A NET873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT874_A NET874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT875_A NET875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT876_A NET876 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT877_A NET877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT878_A NET878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT879_A NET879 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT880_A NET880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT881_A NET881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT882_A NET882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT883_A NET883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT884_A NET884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT885_A NET885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT886_A NET886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT887_A NET887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT888_A NET888 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT889_A NET889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT890_A NET890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT891_A NET891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT892_A NET892 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT893_A NET893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT894_A NET894 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT895_A NET895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT896_A NET896 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT897_A NET897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT898_A NET898 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT899_A NET899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT900_A NET900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT901_A NET901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT902_A NET902 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT903_A NET903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT904_A NET904 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT905_A NET905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT906_A NET906 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT907_A NET907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT908_A NET908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT909_A NET909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT910_A NET910 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT911_A NET911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT912_A NET912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT913_A NET913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT914_A NET914 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT915_A NET915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT916_A NET916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT917_A NET917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT918_A NET918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT919_A NET919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT920_A NET920 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT921_A NET921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT922_A NET922 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT923_A NET923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT924_A NET924 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT925_A NET925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT926_A NET926 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT927_A NET927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT928_A NET928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT929_A NET929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT930_A NET930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT931_A NET931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT932_A NET932 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT933_A NET933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT934_A NET934 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT935_A NET935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT936_A NET936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT937_A NET937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT938_A NET938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT939_A NET939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT940_A NET940 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT941_A NET941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT942_A NET942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT943_A NET943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT944_A NET944 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT945_A NET945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT946_A NET946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT947_A NET947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT948_A NET948 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT949_A NET949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT950_A NET950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT951_A NET951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT952_A NET952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT953_A NET953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT954_A NET954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT955_A NET955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT956_A NET956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT957_A NET957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT958_A NET958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT959_A NET959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT960_A NET960 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT961_A NET961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT962_A NET962 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT963_A NET963 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT964_A NET964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT965_A NET965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT966_A NET966 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT967_A NET967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT968_A NET968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT969_A NET969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT970_A NET970 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT971_A NET971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT972_A NET972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT973_A NET973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT974_A NET974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT975_A NET975 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT976_A NET976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT977_A NET977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT978_A NET978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT979_A NET979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT980_A NET980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT981_A NET981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT982_A NET982 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT983_A NET983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT984_A NET984 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT985_A NET985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT986_A NET986 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT987_A NET987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT988_A NET988 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT989_A NET989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT990_A NET990 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT991_A NET991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT992_A NET992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT993_A NET993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT994_A NET994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT995_A NET995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT996_A NET996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT997_A NET997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT998_A NET998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_OUTPUT999_A NET999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_REPEATER1125_A WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_BUFFERS[0]_A \USER_IRQ_BAR[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_BUFFERS[1]_A \USER_IRQ_BAR[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_BUFFERS[2]_A \USER_IRQ_BAR[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[0]_A NET624 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[0]_B \MPRJ_LOGIC1[458]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[1]_A NET625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[1]_B \MPRJ_LOGIC1[459]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[2]_A NET626 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_ENA_BUF[2]_B \MPRJ_LOGIC1[460]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[0]_A NET621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[0]_B \USER_IRQ_ENABLE[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[1]_A NET622 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[1]_B \USER_IRQ_ENABLE[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[2]_A NET623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_IRQ_GATES[2]_B \USER_IRQ_ENABLE[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[0]_A \LA_DATA_IN_MPRJ_BAR[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[100]_A \LA_DATA_IN_MPRJ_BAR[100]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[101]_A \LA_DATA_IN_MPRJ_BAR[101]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[102]_A \LA_DATA_IN_MPRJ_BAR[102]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[103]_A \LA_DATA_IN_MPRJ_BAR[103]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[104]_A \LA_DATA_IN_MPRJ_BAR[104]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[105]_A \LA_DATA_IN_MPRJ_BAR[105]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[106]_A \LA_DATA_IN_MPRJ_BAR[106]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[107]_A \LA_DATA_IN_MPRJ_BAR[107]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[108]_A \LA_DATA_IN_MPRJ_BAR[108]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[109]_A \LA_DATA_IN_MPRJ_BAR[109]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[10]_A \LA_DATA_IN_MPRJ_BAR[10]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[110]_A \LA_DATA_IN_MPRJ_BAR[110]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[111]_A \LA_DATA_IN_MPRJ_BAR[111]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[112]_A \LA_DATA_IN_MPRJ_BAR[112]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[113]_A \LA_DATA_IN_MPRJ_BAR[113]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[114]_A \LA_DATA_IN_MPRJ_BAR[114]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[115]_A \LA_DATA_IN_MPRJ_BAR[115]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[116]_A \LA_DATA_IN_MPRJ_BAR[116]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[117]_A \LA_DATA_IN_MPRJ_BAR[117]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[118]_A \LA_DATA_IN_MPRJ_BAR[118]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[119]_A \LA_DATA_IN_MPRJ_BAR[119]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[11]_A \LA_DATA_IN_MPRJ_BAR[11]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[120]_A \LA_DATA_IN_MPRJ_BAR[120]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[121]_A \LA_DATA_IN_MPRJ_BAR[121]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[122]_A \LA_DATA_IN_MPRJ_BAR[122]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[123]_A \LA_DATA_IN_MPRJ_BAR[123]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[124]_A \LA_DATA_IN_MPRJ_BAR[124]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[125]_A \LA_DATA_IN_MPRJ_BAR[125]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[126]_A \LA_DATA_IN_MPRJ_BAR[126]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[127]_A \LA_DATA_IN_MPRJ_BAR[127]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[12]_A \LA_DATA_IN_MPRJ_BAR[12]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[13]_A \LA_DATA_IN_MPRJ_BAR[13]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[14]_A \LA_DATA_IN_MPRJ_BAR[14]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[15]_A \LA_DATA_IN_MPRJ_BAR[15]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[16]_A \LA_DATA_IN_MPRJ_BAR[16]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[17]_A \LA_DATA_IN_MPRJ_BAR[17]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[18]_A \LA_DATA_IN_MPRJ_BAR[18]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[19]_A \LA_DATA_IN_MPRJ_BAR[19]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[1]_A \LA_DATA_IN_MPRJ_BAR[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[20]_A \LA_DATA_IN_MPRJ_BAR[20]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[21]_A \LA_DATA_IN_MPRJ_BAR[21]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[22]_A \LA_DATA_IN_MPRJ_BAR[22]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[23]_A \LA_DATA_IN_MPRJ_BAR[23]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[24]_A \LA_DATA_IN_MPRJ_BAR[24]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[25]_A \LA_DATA_IN_MPRJ_BAR[25]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[26]_A \LA_DATA_IN_MPRJ_BAR[26]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[27]_A \LA_DATA_IN_MPRJ_BAR[27]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[28]_A \LA_DATA_IN_MPRJ_BAR[28]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[29]_A \LA_DATA_IN_MPRJ_BAR[29]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[2]_A \LA_DATA_IN_MPRJ_BAR[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[30]_A \LA_DATA_IN_MPRJ_BAR[30]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[31]_A \LA_DATA_IN_MPRJ_BAR[31]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[32]_A \LA_DATA_IN_MPRJ_BAR[32]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[33]_A \LA_DATA_IN_MPRJ_BAR[33]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[34]_A \LA_DATA_IN_MPRJ_BAR[34]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[35]_A \LA_DATA_IN_MPRJ_BAR[35]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[36]_A \LA_DATA_IN_MPRJ_BAR[36]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[37]_A \LA_DATA_IN_MPRJ_BAR[37]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[38]_A \LA_DATA_IN_MPRJ_BAR[38]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[39]_A \LA_DATA_IN_MPRJ_BAR[39]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[3]_A \LA_DATA_IN_MPRJ_BAR[3]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[40]_A \LA_DATA_IN_MPRJ_BAR[40]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[41]_A \LA_DATA_IN_MPRJ_BAR[41]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[42]_A \LA_DATA_IN_MPRJ_BAR[42]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[43]_A \LA_DATA_IN_MPRJ_BAR[43]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[44]_A \LA_DATA_IN_MPRJ_BAR[44]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[45]_A \LA_DATA_IN_MPRJ_BAR[45]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[46]_A \LA_DATA_IN_MPRJ_BAR[46]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[47]_A \LA_DATA_IN_MPRJ_BAR[47]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[48]_A \LA_DATA_IN_MPRJ_BAR[48]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[49]_A \LA_DATA_IN_MPRJ_BAR[49]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[4]_A \LA_DATA_IN_MPRJ_BAR[4]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[50]_A \LA_DATA_IN_MPRJ_BAR[50]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[51]_A \LA_DATA_IN_MPRJ_BAR[51]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[52]_A \LA_DATA_IN_MPRJ_BAR[52]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[53]_A \LA_DATA_IN_MPRJ_BAR[53]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[54]_A \LA_DATA_IN_MPRJ_BAR[54]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[55]_A \LA_DATA_IN_MPRJ_BAR[55]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[56]_A \LA_DATA_IN_MPRJ_BAR[56]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[57]_A \LA_DATA_IN_MPRJ_BAR[57]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[58]_A \LA_DATA_IN_MPRJ_BAR[58]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[59]_A \LA_DATA_IN_MPRJ_BAR[59]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[5]_A \LA_DATA_IN_MPRJ_BAR[5]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[60]_A \LA_DATA_IN_MPRJ_BAR[60]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[61]_A \LA_DATA_IN_MPRJ_BAR[61]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[62]_A \LA_DATA_IN_MPRJ_BAR[62]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[63]_A \LA_DATA_IN_MPRJ_BAR[63]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[64]_A \LA_DATA_IN_MPRJ_BAR[64]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[65]_A \LA_DATA_IN_MPRJ_BAR[65]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[66]_A \LA_DATA_IN_MPRJ_BAR[66]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[67]_A \LA_DATA_IN_MPRJ_BAR[67]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[68]_A \LA_DATA_IN_MPRJ_BAR[68]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[69]_A \LA_DATA_IN_MPRJ_BAR[69]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[6]_A \LA_DATA_IN_MPRJ_BAR[6]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[70]_A \LA_DATA_IN_MPRJ_BAR[70]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[71]_A \LA_DATA_IN_MPRJ_BAR[71]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[72]_A \LA_DATA_IN_MPRJ_BAR[72]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[73]_A \LA_DATA_IN_MPRJ_BAR[73]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[74]_A \LA_DATA_IN_MPRJ_BAR[74]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[75]_A \LA_DATA_IN_MPRJ_BAR[75]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[76]_A \LA_DATA_IN_MPRJ_BAR[76]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[77]_A \LA_DATA_IN_MPRJ_BAR[77]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[78]_A \LA_DATA_IN_MPRJ_BAR[78]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[79]_A \LA_DATA_IN_MPRJ_BAR[79]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[7]_A \LA_DATA_IN_MPRJ_BAR[7]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[80]_A \LA_DATA_IN_MPRJ_BAR[80]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[81]_A \LA_DATA_IN_MPRJ_BAR[81]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[82]_A \LA_DATA_IN_MPRJ_BAR[82]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[83]_A \LA_DATA_IN_MPRJ_BAR[83]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[84]_A \LA_DATA_IN_MPRJ_BAR[84]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[85]_A \LA_DATA_IN_MPRJ_BAR[85]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[86]_A \LA_DATA_IN_MPRJ_BAR[86]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[87]_A \LA_DATA_IN_MPRJ_BAR[87]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[88]_A \LA_DATA_IN_MPRJ_BAR[88]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[89]_A \LA_DATA_IN_MPRJ_BAR[89]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[8]_A \LA_DATA_IN_MPRJ_BAR[8]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[90]_A \LA_DATA_IN_MPRJ_BAR[90]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[91]_A \LA_DATA_IN_MPRJ_BAR[91]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[92]_A \LA_DATA_IN_MPRJ_BAR[92]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[93]_A \LA_DATA_IN_MPRJ_BAR[93]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[94]_A \LA_DATA_IN_MPRJ_BAR[94]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[95]_A \LA_DATA_IN_MPRJ_BAR[95]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[96]_A \LA_DATA_IN_MPRJ_BAR[96]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[97]_A \LA_DATA_IN_MPRJ_BAR[97]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[98]_A \LA_DATA_IN_MPRJ_BAR[98]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[99]_A \LA_DATA_IN_MPRJ_BAR[99]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_BUFFERS[9]_A \LA_DATA_IN_MPRJ_BAR[9]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[0]_A NET260 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[0]_B \MPRJ_LOGIC1[330]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[100]_A NET261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[100]_B \MPRJ_LOGIC1[430]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[101]_A NET262 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[101]_B \MPRJ_LOGIC1[431]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[102]_A NET263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[102]_B \MPRJ_LOGIC1[432]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[103]_A NET264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[103]_B \MPRJ_LOGIC1[433]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[104]_A NET265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[104]_B \MPRJ_LOGIC1[434]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[105]_A NET266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[105]_B \MPRJ_LOGIC1[435]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[106]_A NET267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[106]_B \MPRJ_LOGIC1[436]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[107]_A NET268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[107]_B \MPRJ_LOGIC1[437]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[108]_A NET269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[108]_B \MPRJ_LOGIC1[438]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[109]_A NET270 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[109]_B \MPRJ_LOGIC1[439]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[10]_A NET271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[10]_B \MPRJ_LOGIC1[340]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[110]_A NET272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[110]_B \MPRJ_LOGIC1[440]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[111]_A NET273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[111]_B \MPRJ_LOGIC1[441]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[112]_A NET274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[112]_B \MPRJ_LOGIC1[442]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[113]_A NET275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[113]_B \MPRJ_LOGIC1[443]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[114]_A NET276 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[114]_B \MPRJ_LOGIC1[444]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[115]_A NET277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[115]_B \MPRJ_LOGIC1[445]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[116]_A NET278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[116]_B \MPRJ_LOGIC1[446]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[117]_A NET279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[117]_B \MPRJ_LOGIC1[447]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[118]_A NET280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[118]_B \MPRJ_LOGIC1[448]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[119]_A NET281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[119]_B \MPRJ_LOGIC1[449]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[11]_A NET282 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[11]_B \MPRJ_LOGIC1[341]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[120]_A NET283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[120]_B \MPRJ_LOGIC1[450]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[121]_A NET284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[121]_B \MPRJ_LOGIC1[451]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[122]_A NET285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[122]_B \MPRJ_LOGIC1[452]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[123]_A NET286 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[123]_B \MPRJ_LOGIC1[453]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[124]_A NET287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[124]_B \MPRJ_LOGIC1[454]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[125]_A NET288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[125]_B \MPRJ_LOGIC1[455]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[126]_A NET289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[126]_B \MPRJ_LOGIC1[456]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[127]_A NET290 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[127]_B \MPRJ_LOGIC1[457]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[12]_A NET291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[12]_B \MPRJ_LOGIC1[342]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[13]_A NET292 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[13]_B \MPRJ_LOGIC1[343]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[14]_A NET293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[14]_B \MPRJ_LOGIC1[344]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[15]_A NET294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[15]_B \MPRJ_LOGIC1[345]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[16]_A NET295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[16]_B \MPRJ_LOGIC1[346]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[17]_A NET296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[17]_B \MPRJ_LOGIC1[347]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[18]_A NET297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[18]_B \MPRJ_LOGIC1[348]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[19]_A NET298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[19]_B \MPRJ_LOGIC1[349]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[1]_A NET299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[1]_B \MPRJ_LOGIC1[331]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[20]_A NET300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[20]_B \MPRJ_LOGIC1[350]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[21]_A NET301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[21]_B \MPRJ_LOGIC1[351]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[22]_A NET302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[22]_B \MPRJ_LOGIC1[352]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[23]_A NET303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[23]_B \MPRJ_LOGIC1[353]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[24]_A NET304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[24]_B \MPRJ_LOGIC1[354]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[25]_A NET305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[25]_B \MPRJ_LOGIC1[355]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[26]_A NET306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[26]_B \MPRJ_LOGIC1[356]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[27]_A NET307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[27]_B \MPRJ_LOGIC1[357]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[28]_A NET308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[28]_B \MPRJ_LOGIC1[358]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[29]_A NET309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[29]_B \MPRJ_LOGIC1[359]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[2]_A NET310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[2]_B \MPRJ_LOGIC1[332]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[30]_A NET311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[30]_B \MPRJ_LOGIC1[360]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[31]_A NET312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[31]_B \MPRJ_LOGIC1[361]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[32]_A NET313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[32]_B \MPRJ_LOGIC1[362]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[33]_A NET314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[33]_B \MPRJ_LOGIC1[363]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[34]_A NET315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[34]_B \MPRJ_LOGIC1[364]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[35]_A NET316 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[35]_B \MPRJ_LOGIC1[365]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[36]_A NET317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[36]_B \MPRJ_LOGIC1[366]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[37]_A NET318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[37]_B \MPRJ_LOGIC1[367]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[38]_A NET319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[38]_B \MPRJ_LOGIC1[368]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[39]_A NET320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[39]_B \MPRJ_LOGIC1[369]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[3]_A NET321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[3]_B \MPRJ_LOGIC1[333]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[40]_A NET322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[40]_B \MPRJ_LOGIC1[370]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[41]_A NET323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[41]_B \MPRJ_LOGIC1[371]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[42]_A NET324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[42]_B \MPRJ_LOGIC1[372]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[43]_A NET325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[43]_B \MPRJ_LOGIC1[373]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[44]_A NET326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[44]_B \MPRJ_LOGIC1[374]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[45]_A NET327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[45]_B \MPRJ_LOGIC1[375]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[46]_A NET328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[46]_B \MPRJ_LOGIC1[376]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[47]_A NET329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[47]_B \MPRJ_LOGIC1[377]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[48]_A NET330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[48]_B \MPRJ_LOGIC1[378]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[49]_A NET331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[49]_B \MPRJ_LOGIC1[379]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[4]_A NET332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[4]_B \MPRJ_LOGIC1[334]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[50]_A NET333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[50]_B \MPRJ_LOGIC1[380]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[51]_A NET334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[51]_B \MPRJ_LOGIC1[381]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[52]_A NET335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[52]_B \MPRJ_LOGIC1[382]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[53]_A NET336 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[53]_B \MPRJ_LOGIC1[383]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[54]_A NET337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[54]_B \MPRJ_LOGIC1[384]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[55]_A NET338 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[55]_B \MPRJ_LOGIC1[385]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[56]_A NET339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[56]_B \MPRJ_LOGIC1[386]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[57]_A NET340 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[57]_B \MPRJ_LOGIC1[387]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[58]_A NET341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[58]_B \MPRJ_LOGIC1[388]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[59]_A NET342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[59]_B \MPRJ_LOGIC1[389]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[5]_A NET343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[5]_B \MPRJ_LOGIC1[335]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[60]_A NET344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[60]_B \MPRJ_LOGIC1[390]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[61]_A NET345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[61]_B \MPRJ_LOGIC1[391]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[62]_A NET346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[62]_B \MPRJ_LOGIC1[392]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[63]_A NET347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[63]_B \MPRJ_LOGIC1[393]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[64]_A NET348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[64]_B \MPRJ_LOGIC1[394]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[65]_A NET349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[65]_B \MPRJ_LOGIC1[395]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[66]_A NET350 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[66]_B \MPRJ_LOGIC1[396]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[67]_A NET351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[67]_B \MPRJ_LOGIC1[397]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[68]_A NET352 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[68]_B \MPRJ_LOGIC1[398]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[69]_A NET353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[69]_B \MPRJ_LOGIC1[399]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[6]_A NET354 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[6]_B \MPRJ_LOGIC1[336]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[70]_A NET355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[70]_B \MPRJ_LOGIC1[400]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[71]_A NET356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[71]_B \MPRJ_LOGIC1[401]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[72]_A NET357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[72]_B \MPRJ_LOGIC1[402]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[73]_A NET358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[73]_B \MPRJ_LOGIC1[403]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[74]_A NET359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[74]_B \MPRJ_LOGIC1[404]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[75]_A NET360 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[75]_B \MPRJ_LOGIC1[405]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[76]_A NET361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[76]_B \MPRJ_LOGIC1[406]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[77]_A NET362 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[77]_B \MPRJ_LOGIC1[407]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[78]_A NET363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[78]_B \MPRJ_LOGIC1[408]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[79]_A NET364 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[79]_B \MPRJ_LOGIC1[409]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[7]_A NET365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[7]_B \MPRJ_LOGIC1[337]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[80]_A NET366 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[80]_B \MPRJ_LOGIC1[410]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[81]_A NET367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[81]_B \MPRJ_LOGIC1[411]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[82]_A NET368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[82]_B \MPRJ_LOGIC1[412]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[83]_A NET369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[83]_B \MPRJ_LOGIC1[413]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[84]_A NET370 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[84]_B \MPRJ_LOGIC1[414]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[85]_A NET371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[85]_B \MPRJ_LOGIC1[415]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[86]_A NET372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[86]_B \MPRJ_LOGIC1[416]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[87]_A NET373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[87]_B \MPRJ_LOGIC1[417]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[88]_A NET374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[88]_B \MPRJ_LOGIC1[418]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[89]_A NET375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[89]_B \MPRJ_LOGIC1[419]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[8]_A NET376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[8]_B \MPRJ_LOGIC1[338]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[90]_A NET377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[90]_B \MPRJ_LOGIC1[420]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[91]_A NET378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[91]_B \MPRJ_LOGIC1[421]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[92]_A NET379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[92]_B \MPRJ_LOGIC1[422]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[93]_A NET380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[93]_B \MPRJ_LOGIC1[423]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[94]_A NET381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[94]_B \MPRJ_LOGIC1[424]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[95]_A NET382 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[95]_B \MPRJ_LOGIC1[425]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[96]_A NET383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[96]_B \MPRJ_LOGIC1[426]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[97]_A NET384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[97]_B \MPRJ_LOGIC1[427]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[98]_A NET385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[98]_B \MPRJ_LOGIC1[428]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[99]_A NET386 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[99]_B \MPRJ_LOGIC1[429]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[9]_A NET387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_ENA_BUF[9]_B \MPRJ_LOGIC1[339]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[0]_A NET4 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[0]_B \LA_DATA_IN_ENABLE[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[100]_A NET5 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[100]_B \LA_DATA_IN_ENABLE[100]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[101]_A NET6 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[101]_B \LA_DATA_IN_ENABLE[101]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[102]_A NET7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[102]_B \LA_DATA_IN_ENABLE[102]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[103]_A NET8 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[103]_B \LA_DATA_IN_ENABLE[103]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[104]_A NET9 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[104]_B \LA_DATA_IN_ENABLE[104]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[105]_A NET10 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[105]_B \LA_DATA_IN_ENABLE[105]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[106]_A NET11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[106]_B \LA_DATA_IN_ENABLE[106]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[107]_A NET12 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[107]_B \LA_DATA_IN_ENABLE[107]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[108]_A NET13 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[108]_B \LA_DATA_IN_ENABLE[108]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[109]_A NET14 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[109]_B \LA_DATA_IN_ENABLE[109]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[10]_A NET15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[10]_B \LA_DATA_IN_ENABLE[10]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[110]_A NET16 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[110]_B \LA_DATA_IN_ENABLE[110]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[111]_A NET17 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[111]_B \LA_DATA_IN_ENABLE[111]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[112]_A NET18 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[112]_B \LA_DATA_IN_ENABLE[112]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[113]_A NET19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[113]_B \LA_DATA_IN_ENABLE[113]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[114]_A NET20 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[114]_B \LA_DATA_IN_ENABLE[114]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[115]_A NET21 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[115]_B \LA_DATA_IN_ENABLE[115]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[116]_A NET22 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[116]_B \LA_DATA_IN_ENABLE[116]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[117]_A NET23 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[117]_B \LA_DATA_IN_ENABLE[117]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[118]_A NET24 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[118]_B \LA_DATA_IN_ENABLE[118]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[119]_A NET25 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[119]_B \LA_DATA_IN_ENABLE[119]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[11]_A NET26 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[11]_B \LA_DATA_IN_ENABLE[11]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[120]_A NET27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[120]_B \LA_DATA_IN_ENABLE[120]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[121]_A NET28 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[121]_B \LA_DATA_IN_ENABLE[121]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[122]_A NET29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[122]_B \LA_DATA_IN_ENABLE[122]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[123]_A NET30 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[123]_B \LA_DATA_IN_ENABLE[123]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[124]_A NET31 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[124]_B \LA_DATA_IN_ENABLE[124]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[125]_A NET32 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[125]_B \LA_DATA_IN_ENABLE[125]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[126]_A NET33 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[126]_B \LA_DATA_IN_ENABLE[126]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[127]_A NET34 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[127]_B \LA_DATA_IN_ENABLE[127]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[12]_A NET35 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[12]_B \LA_DATA_IN_ENABLE[12]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[13]_A NET36 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[13]_B \LA_DATA_IN_ENABLE[13]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[14]_A NET37 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[14]_B \LA_DATA_IN_ENABLE[14]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[15]_A NET38 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[15]_B \LA_DATA_IN_ENABLE[15]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[16]_A NET39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[16]_B \LA_DATA_IN_ENABLE[16]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[17]_A NET40 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[17]_B \LA_DATA_IN_ENABLE[17]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[18]_A NET41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[18]_B \LA_DATA_IN_ENABLE[18]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[19]_A NET42 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[19]_B \LA_DATA_IN_ENABLE[19]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[1]_A NET43 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[1]_B \LA_DATA_IN_ENABLE[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[20]_A NET44 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[20]_B \LA_DATA_IN_ENABLE[20]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[21]_A NET45 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[21]_B \LA_DATA_IN_ENABLE[21]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[22]_A NET46 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[22]_B \LA_DATA_IN_ENABLE[22]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[23]_A NET47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[23]_B \LA_DATA_IN_ENABLE[23]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[24]_A NET48 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[24]_B \LA_DATA_IN_ENABLE[24]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[25]_A NET49 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[25]_B \LA_DATA_IN_ENABLE[25]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[26]_A NET50 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[26]_B \LA_DATA_IN_ENABLE[26]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[27]_A NET51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[27]_B \LA_DATA_IN_ENABLE[27]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[28]_A NET52 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[28]_B \LA_DATA_IN_ENABLE[28]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[29]_A NET53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[29]_B \LA_DATA_IN_ENABLE[29]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[2]_A NET54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[2]_B \LA_DATA_IN_ENABLE[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[30]_A NET55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[30]_B \LA_DATA_IN_ENABLE[30]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[31]_A NET56 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[31]_B \LA_DATA_IN_ENABLE[31]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[32]_A NET57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[32]_B \LA_DATA_IN_ENABLE[32]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[33]_A NET58 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[33]_B \LA_DATA_IN_ENABLE[33]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[34]_A NET59 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[34]_B \LA_DATA_IN_ENABLE[34]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[35]_A NET60 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[35]_B \LA_DATA_IN_ENABLE[35]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[36]_A NET61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[36]_B \LA_DATA_IN_ENABLE[36]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[37]_A NET62 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[37]_B \LA_DATA_IN_ENABLE[37]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[38]_A NET63 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[38]_B \LA_DATA_IN_ENABLE[38]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[39]_A NET64 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[39]_B \LA_DATA_IN_ENABLE[39]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[3]_A NET65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[3]_B \LA_DATA_IN_ENABLE[3]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[40]_A NET66 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[40]_B \LA_DATA_IN_ENABLE[40]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[41]_A NET67 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[41]_B \LA_DATA_IN_ENABLE[41]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[42]_A NET68 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[42]_B \LA_DATA_IN_ENABLE[42]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[43]_A NET69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[43]_B \LA_DATA_IN_ENABLE[43]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[44]_A NET70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[44]_B \LA_DATA_IN_ENABLE[44]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[45]_A NET71 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[45]_B \LA_DATA_IN_ENABLE[45]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[46]_A NET72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[46]_B \LA_DATA_IN_ENABLE[46]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[47]_A NET73 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[47]_B \LA_DATA_IN_ENABLE[47]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[48]_A NET74 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[48]_B \LA_DATA_IN_ENABLE[48]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[49]_A NET75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[49]_B \LA_DATA_IN_ENABLE[49]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[4]_A NET76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[4]_B \LA_DATA_IN_ENABLE[4]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[50]_A NET77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[50]_B \LA_DATA_IN_ENABLE[50]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[51]_A NET78 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[51]_B \LA_DATA_IN_ENABLE[51]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[52]_A NET79 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[52]_B \LA_DATA_IN_ENABLE[52]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[53]_A NET80 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[53]_B \LA_DATA_IN_ENABLE[53]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[54]_A NET81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[54]_B \LA_DATA_IN_ENABLE[54]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[55]_A NET82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[55]_B \LA_DATA_IN_ENABLE[55]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[56]_A NET83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[56]_B \LA_DATA_IN_ENABLE[56]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[57]_A NET84 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[57]_B \LA_DATA_IN_ENABLE[57]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[58]_A NET85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[58]_B \LA_DATA_IN_ENABLE[58]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[59]_A NET86 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[59]_B \LA_DATA_IN_ENABLE[59]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[5]_A NET87 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[5]_B \LA_DATA_IN_ENABLE[5]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[60]_A NET88 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[60]_B \LA_DATA_IN_ENABLE[60]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[61]_A NET89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[61]_B \LA_DATA_IN_ENABLE[61]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[62]_A NET90 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[62]_B \LA_DATA_IN_ENABLE[62]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[63]_A NET91 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[63]_B \LA_DATA_IN_ENABLE[63]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[64]_A NET92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[64]_B \LA_DATA_IN_ENABLE[64]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[65]_A NET93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[65]_B \LA_DATA_IN_ENABLE[65]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[66]_A NET94 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[66]_B \LA_DATA_IN_ENABLE[66]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[67]_A NET95 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[67]_B \LA_DATA_IN_ENABLE[67]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[68]_A NET96 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[68]_B \LA_DATA_IN_ENABLE[68]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[69]_A NET97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[69]_B \LA_DATA_IN_ENABLE[69]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[6]_A NET98 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[6]_B \LA_DATA_IN_ENABLE[6]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[70]_A NET99 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[70]_B \LA_DATA_IN_ENABLE[70]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[71]_A NET100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[71]_B \LA_DATA_IN_ENABLE[71]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[72]_A NET101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[72]_B \LA_DATA_IN_ENABLE[72]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[73]_A NET102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[73]_B \LA_DATA_IN_ENABLE[73]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[74]_A NET103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[74]_B \LA_DATA_IN_ENABLE[74]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[75]_A NET104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[75]_B \LA_DATA_IN_ENABLE[75]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[76]_A NET105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[76]_B \LA_DATA_IN_ENABLE[76]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[77]_A NET106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[77]_B \LA_DATA_IN_ENABLE[77]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[78]_A NET107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[78]_B \LA_DATA_IN_ENABLE[78]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[79]_A NET108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[79]_B \LA_DATA_IN_ENABLE[79]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[7]_A NET109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[7]_B \LA_DATA_IN_ENABLE[7]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[80]_A NET110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[80]_B \LA_DATA_IN_ENABLE[80]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[81]_A NET111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[81]_B \LA_DATA_IN_ENABLE[81]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[82]_A NET112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[82]_B \LA_DATA_IN_ENABLE[82]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[83]_A NET113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[83]_B \LA_DATA_IN_ENABLE[83]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[84]_A NET114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[84]_B \LA_DATA_IN_ENABLE[84]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[85]_A NET115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[85]_B \LA_DATA_IN_ENABLE[85]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[86]_A NET116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[86]_B \LA_DATA_IN_ENABLE[86]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[87]_A NET117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[87]_B \LA_DATA_IN_ENABLE[87]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[88]_A NET118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[88]_B \LA_DATA_IN_ENABLE[88]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[89]_A NET119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[89]_B \LA_DATA_IN_ENABLE[89]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[8]_A NET120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[8]_B \LA_DATA_IN_ENABLE[8]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[90]_A NET121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[90]_B \LA_DATA_IN_ENABLE[90]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[91]_A NET122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[91]_B \LA_DATA_IN_ENABLE[91]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[92]_A NET123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[92]_B \LA_DATA_IN_ENABLE[92]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[93]_A NET124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[93]_B \LA_DATA_IN_ENABLE[93]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[94]_A NET125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[94]_B \LA_DATA_IN_ENABLE[94]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[95]_A NET126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[95]_B \LA_DATA_IN_ENABLE[95]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[96]_A NET127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[96]_B \LA_DATA_IN_ENABLE[96]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[97]_A NET128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[97]_B \LA_DATA_IN_ENABLE[97]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[98]_A NET129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[98]_B \LA_DATA_IN_ENABLE[98]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[99]_A NET130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[99]_B \LA_DATA_IN_ENABLE[99]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[9]_A NET131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_IN_GATES[9]_B \LA_DATA_IN_ENABLE[9]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[0]_A _201_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[0]_TE \MPRJ_LOGIC1[202]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[100]_A _202_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[100]_TE \MPRJ_LOGIC1[302]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[101]_A _203_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[101]_TE \MPRJ_LOGIC1[303]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[102]_A _204_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[102]_TE \MPRJ_LOGIC1[304]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[103]_A _205_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[103]_TE \MPRJ_LOGIC1[305]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[104]_A _206_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[104]_TE \MPRJ_LOGIC1[306]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[105]_A _207_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[105]_TE \MPRJ_LOGIC1[307]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[106]_A _208_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[106]_TE \MPRJ_LOGIC1[308]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[107]_A _209_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[107]_TE \MPRJ_LOGIC1[309]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[108]_A _210_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[108]_TE \MPRJ_LOGIC1[310]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[109]_A _211_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[109]_TE \MPRJ_LOGIC1[311]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[10]_A _212_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[10]_TE \MPRJ_LOGIC1[212]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[110]_A _213_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[110]_TE \MPRJ_LOGIC1[312]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[111]_A _214_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[111]_TE \MPRJ_LOGIC1[313]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[112]_A _215_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[112]_TE \MPRJ_LOGIC1[314]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[113]_A _216_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[113]_TE \MPRJ_LOGIC1[315]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[114]_A _217_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[114]_TE \MPRJ_LOGIC1[316]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[115]_A _218_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[115]_TE \MPRJ_LOGIC1[317]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[116]_A _219_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[116]_TE \MPRJ_LOGIC1[318]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[117]_A _220_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[117]_TE \MPRJ_LOGIC1[319]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[118]_A _221_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[118]_TE \MPRJ_LOGIC1[320]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[119]_A _222_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[119]_TE \MPRJ_LOGIC1[321]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[11]_A _223_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[11]_TE \MPRJ_LOGIC1[213]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[120]_A _224_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[120]_TE \MPRJ_LOGIC1[322]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[121]_A _225_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[121]_TE \MPRJ_LOGIC1[323]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[122]_A _226_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[122]_TE \MPRJ_LOGIC1[324]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[123]_A _227_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[123]_TE \MPRJ_LOGIC1[325]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[124]_A _228_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[124]_TE \MPRJ_LOGIC1[326]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[125]_A _229_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[125]_TE \MPRJ_LOGIC1[327]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[126]_A _230_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[126]_TE \MPRJ_LOGIC1[328]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[127]_A _231_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[127]_TE \MPRJ_LOGIC1[329]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[12]_A _232_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[12]_TE \MPRJ_LOGIC1[214]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[13]_A _233_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[13]_TE \MPRJ_LOGIC1[215]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[14]_A _234_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[14]_TE \MPRJ_LOGIC1[216]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[15]_A _235_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[15]_TE \MPRJ_LOGIC1[217]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[16]_A _236_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[16]_TE \MPRJ_LOGIC1[218]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[17]_A _237_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[17]_TE \MPRJ_LOGIC1[219]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[18]_A _238_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[18]_TE \MPRJ_LOGIC1[220]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[19]_A _239_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[19]_TE \MPRJ_LOGIC1[221]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[1]_A _240_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[1]_TE \MPRJ_LOGIC1[203]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[20]_A _241_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[20]_TE \MPRJ_LOGIC1[222]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[21]_A _242_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[21]_TE \MPRJ_LOGIC1[223]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[22]_A _243_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[22]_TE \MPRJ_LOGIC1[224]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[23]_A _244_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[23]_TE \MPRJ_LOGIC1[225]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[24]_A _245_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[24]_TE \MPRJ_LOGIC1[226]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[25]_A _246_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[25]_TE \MPRJ_LOGIC1[227]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[26]_A _247_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[26]_TE \MPRJ_LOGIC1[228]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[27]_A _248_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[27]_TE \MPRJ_LOGIC1[229]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[28]_A _249_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[28]_TE \MPRJ_LOGIC1[230]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[29]_A _250_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[29]_TE \MPRJ_LOGIC1[231]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[2]_A _251_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[2]_TE \MPRJ_LOGIC1[204]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[30]_A _252_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[30]_TE \MPRJ_LOGIC1[232]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[31]_A _253_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[31]_TE \MPRJ_LOGIC1[233]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[32]_A _254_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[32]_TE \MPRJ_LOGIC1[234]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[33]_A _255_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[33]_TE \MPRJ_LOGIC1[235]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[34]_A _256_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[34]_TE \MPRJ_LOGIC1[236]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[35]_A _257_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[35]_TE \MPRJ_LOGIC1[237]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[36]_A _258_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[36]_TE \MPRJ_LOGIC1[238]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[37]_A _259_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[37]_TE \MPRJ_LOGIC1[239]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[38]_A _260_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[38]_TE \MPRJ_LOGIC1[240]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[39]_A _261_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[39]_TE \MPRJ_LOGIC1[241]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[3]_A _262_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[3]_TE \MPRJ_LOGIC1[205]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[40]_A _263_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[40]_TE \MPRJ_LOGIC1[242]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[41]_A _264_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[41]_TE \MPRJ_LOGIC1[243]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[42]_A _265_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[42]_TE \MPRJ_LOGIC1[244]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[43]_A _266_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[43]_TE \MPRJ_LOGIC1[245]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[44]_A _267_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[44]_TE \MPRJ_LOGIC1[246]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[45]_A _268_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[45]_TE \MPRJ_LOGIC1[247]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[46]_A _269_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[46]_TE \MPRJ_LOGIC1[248]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[47]_A _270_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[47]_TE \MPRJ_LOGIC1[249]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[48]_A _271_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[48]_TE \MPRJ_LOGIC1[250]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[49]_A _272_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[49]_TE \MPRJ_LOGIC1[251]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[4]_A _273_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[4]_TE \MPRJ_LOGIC1[206]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[50]_A _274_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[50]_TE \MPRJ_LOGIC1[252]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[51]_A _275_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[51]_TE \MPRJ_LOGIC1[253]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[52]_A _276_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[52]_TE \MPRJ_LOGIC1[254]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[53]_A _277_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[53]_TE \MPRJ_LOGIC1[255]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[54]_A _278_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[54]_TE \MPRJ_LOGIC1[256]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[55]_A _279_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[55]_TE \MPRJ_LOGIC1[257]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[56]_A _280_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[56]_TE \MPRJ_LOGIC1[258]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[57]_A _281_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[57]_TE \MPRJ_LOGIC1[259]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[58]_A _282_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[58]_TE \MPRJ_LOGIC1[260]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[59]_A _283_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[59]_TE \MPRJ_LOGIC1[261]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[5]_A _284_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[5]_TE \MPRJ_LOGIC1[207]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[60]_A _285_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[60]_TE \MPRJ_LOGIC1[262]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[61]_A _286_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[61]_TE \MPRJ_LOGIC1[263]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[62]_A _287_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[62]_TE \MPRJ_LOGIC1[264]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[63]_A _288_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[63]_TE \MPRJ_LOGIC1[265]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[64]_A _289_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[64]_TE \MPRJ_LOGIC1[266]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[65]_A _290_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[65]_TE \MPRJ_LOGIC1[267]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[66]_A _291_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[66]_TE \MPRJ_LOGIC1[268]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[67]_A _292_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[67]_TE \MPRJ_LOGIC1[269]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[68]_A _293_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[68]_TE \MPRJ_LOGIC1[270]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[69]_A _294_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[69]_TE \MPRJ_LOGIC1[271]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[6]_A _295_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[6]_TE \MPRJ_LOGIC1[208]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[70]_A _296_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[70]_TE \MPRJ_LOGIC1[272]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[71]_A _297_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[71]_TE \MPRJ_LOGIC1[273]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[72]_A _298_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[72]_TE \MPRJ_LOGIC1[274]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[73]_A _299_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[73]_TE \MPRJ_LOGIC1[275]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[74]_A _300_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[74]_TE \MPRJ_LOGIC1[276]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[75]_A _301_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[75]_TE \MPRJ_LOGIC1[277]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[76]_A _302_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[76]_TE \MPRJ_LOGIC1[278]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[77]_A _303_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[77]_TE \MPRJ_LOGIC1[279]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[78]_A _304_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[78]_TE \MPRJ_LOGIC1[280]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[79]_A _305_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[79]_TE \MPRJ_LOGIC1[281]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[7]_A _306_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[7]_TE \MPRJ_LOGIC1[209]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[80]_A _307_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[80]_TE \MPRJ_LOGIC1[282]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[81]_A _308_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[81]_TE \MPRJ_LOGIC1[283]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[82]_A _309_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[82]_TE \MPRJ_LOGIC1[284]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[83]_A _310_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[83]_TE \MPRJ_LOGIC1[285]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[84]_A _311_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[84]_TE \MPRJ_LOGIC1[286]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[85]_A _312_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[85]_TE \MPRJ_LOGIC1[287]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[86]_A _313_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[86]_TE \MPRJ_LOGIC1[288]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[87]_A _314_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[87]_TE \MPRJ_LOGIC1[289]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[88]_A _315_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[88]_TE \MPRJ_LOGIC1[290]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[89]_A _316_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[89]_TE \MPRJ_LOGIC1[291]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[8]_A _317_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[8]_TE \MPRJ_LOGIC1[210]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[90]_A _318_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[90]_TE \MPRJ_LOGIC1[292]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[91]_A _319_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[91]_TE \MPRJ_LOGIC1[293]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[92]_A _320_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[92]_TE \MPRJ_LOGIC1[294]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[93]_A _321_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[93]_TE \MPRJ_LOGIC1[295]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[94]_A _322_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[94]_TE \MPRJ_LOGIC1[296]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[95]_A _323_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[95]_TE \MPRJ_LOGIC1[297]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[96]_A _324_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[96]_TE \MPRJ_LOGIC1[298]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[97]_A _325_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[97]_TE \MPRJ_LOGIC1[299]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[98]_A _326_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[98]_TE \MPRJ_LOGIC1[300]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[99]_A _327_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[99]_TE \MPRJ_LOGIC1[301]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[9]_A _328_ VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_TO_MPRJ_OEN_BUFFERS[9]_TE \MPRJ_LOGIC1[211]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_USER_TO_MPRJ_WB_ENA_BUF_A NET614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_USER_TO_MPRJ_WB_ENA_BUF_B \MPRJ_LOGIC1[462]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_USER_WB_ACK_BUFFER_A MPRJ_ACK_I_CORE_BAR VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_USER_WB_ACK_GATE_A NET516 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XANTENNA_USER_WB_ACK_GATE_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[0]_A \MPRJ_DAT_I_CORE_BAR[0]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[10]_A \MPRJ_DAT_I_CORE_BAR[10]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[11]_A \MPRJ_DAT_I_CORE_BAR[11]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[12]_A \MPRJ_DAT_I_CORE_BAR[12]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[13]_A \MPRJ_DAT_I_CORE_BAR[13]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[14]_A \MPRJ_DAT_I_CORE_BAR[14]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[15]_A \MPRJ_DAT_I_CORE_BAR[15]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[16]_A \MPRJ_DAT_I_CORE_BAR[16]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[17]_A \MPRJ_DAT_I_CORE_BAR[17]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[18]_A \MPRJ_DAT_I_CORE_BAR[18]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[19]_A \MPRJ_DAT_I_CORE_BAR[19]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[1]_A \MPRJ_DAT_I_CORE_BAR[1]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[20]_A \MPRJ_DAT_I_CORE_BAR[20]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[21]_A \MPRJ_DAT_I_CORE_BAR[21]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[22]_A \MPRJ_DAT_I_CORE_BAR[22]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[23]_A \MPRJ_DAT_I_CORE_BAR[23]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[24]_A \MPRJ_DAT_I_CORE_BAR[24]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[25]_A \MPRJ_DAT_I_CORE_BAR[25]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[26]_A \MPRJ_DAT_I_CORE_BAR[26]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[27]_A \MPRJ_DAT_I_CORE_BAR[27]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[28]_A \MPRJ_DAT_I_CORE_BAR[28]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[29]_A \MPRJ_DAT_I_CORE_BAR[29]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[2]_A \MPRJ_DAT_I_CORE_BAR[2]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[30]_A \MPRJ_DAT_I_CORE_BAR[30]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[31]_A \MPRJ_DAT_I_CORE_BAR[31]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[3]_A \MPRJ_DAT_I_CORE_BAR[3]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[4]_A \MPRJ_DAT_I_CORE_BAR[4]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[5]_A \MPRJ_DAT_I_CORE_BAR[5]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[6]_A \MPRJ_DAT_I_CORE_BAR[6]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[7]_A \MPRJ_DAT_I_CORE_BAR[7]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[8]_A \MPRJ_DAT_I_CORE_BAR[8]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_BUFFERS[9]_A \MPRJ_DAT_I_CORE_BAR[9]  VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[0]_A NET550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[0]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[10]_A NET551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[10]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[11]_A NET552 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[11]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[12]_A NET553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[12]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[13]_A NET554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[13]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[14]_A NET555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[14]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[15]_A NET556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[15]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[16]_A NET557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[16]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[17]_A NET558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[17]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[18]_A NET559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[18]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[19]_A NET560 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[19]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[1]_A NET561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[1]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[20]_A NET562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[20]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[21]_A NET563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[21]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[22]_A NET564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[22]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[23]_A NET565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[23]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[24]_A NET566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[24]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[25]_A NET567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[25]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[26]_A NET568 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[26]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[27]_A NET569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[27]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[28]_A NET570 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[28]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[29]_A NET571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[29]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[2]_A NET572 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[2]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[30]_A NET573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[30]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[31]_A NET574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[31]_B NET1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[3]_A NET575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[3]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[4]_A NET576 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[4]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[5]_A NET577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[5]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[6]_A NET578 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[6]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[7]_A NET579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[7]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[8]_A NET580 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[8]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[9]_A NET581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
X\ANTENNA_USER_WB_DAT_GATES[9]_B WB_IN_ENABLE VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DIODE_2
XFILLER_0_1030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1224 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1270 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1286 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1534 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1580 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1728 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2042 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2142 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2290 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_0_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_2346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_240 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_736 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_0_946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_0_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_10_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1047 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_10_1115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1386 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1446 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1535 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1610 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_10_1835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_400 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_404 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_428 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_10_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_846 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_850 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_858 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_862 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_10_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_10_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_10_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_10_957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_10_969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_10_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1046 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_11_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_11_1489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_1508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_1850 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_1858 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1870 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_514 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_11_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_11_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_11_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_11_817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_844 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_11_854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_11_972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_11_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_11_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1602 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_1606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1630 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_12_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_12_1702 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_1706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_1710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_12_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_12_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_12_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_12_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_12_579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_12_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_12_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_12_656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_12_664 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_12_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_12_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_12_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_13_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_13_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_13_1723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_13_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1879 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_13_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_1975 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_13_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_13_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_13_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_13_632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_636 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_13_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_13_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_13_655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_13_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_13_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_13_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_14_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_1616 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_14_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_14_1687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_14_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_1732 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1736 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_14_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_14_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_14_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_14_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_1975 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_14_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_14_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_14_668 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_14_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_14_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_14_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_14_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_1556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1560 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1576 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1600 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_15_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_15_1710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1714 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_15_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_1879 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_15_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_2005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_2008 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_15_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_15_519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_15_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_15_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_599 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_15_639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_15_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_652 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_15_656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_668 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_680 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_15_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_15_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_15_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_15_730 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_16_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1600 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_16_1699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_16_1740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_16_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_16_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_16_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1888 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_1904 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_1940 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1944 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_16_530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_534 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_16_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_16_647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_16_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_16_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_16_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_16_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_17_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_17_1639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_17_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_17_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1750 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1766 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_17_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_17_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_17_563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_17_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_17_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_17_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_17_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_17_654 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_17_662 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_686 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_17_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_17_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_18_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1598 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1602 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1626 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_18_1724 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1738 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_18_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1896 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1963 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_2003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_18_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_420 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_570 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_594 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_18_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_18_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_18_687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_18_705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_18_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_18_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_18_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1932 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_19_194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1948 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_19_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_19_481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_19_528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_546 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_19_558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_19_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_19_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_19_676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_680 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_19_684 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_696 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_19_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_19_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_19_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_19_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_1_1004 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1014 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1019 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1028 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1047 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1058 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1150 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1438 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1504 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1520 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1535 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1590 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_16 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1612 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1616 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1652 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1678 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1712 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1730 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1784 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1830 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1842 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1864 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1914 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1922 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1926 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_20 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_204 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2082 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2086 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2140 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2214 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_2245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_2350 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_26 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_350 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_36 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_40 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_43 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_476 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_516 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_570 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_578 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_624 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_636 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_686 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_71 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_732 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_818 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_862 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_870 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_888 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_892 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_1_904 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_934 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_1_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_984 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_988 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_1_995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_1_999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_1613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_1783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1786 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_1798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1842 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_20_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_1874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1898 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1910 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_20_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1924 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_1936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1960 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_1977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_232 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_236 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_20_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_20_482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_20_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_20_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_578 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_58 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_20_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_20_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_20_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_20_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_20_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_21_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_140 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_1699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_1742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1746 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1758 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_176 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_1779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1786 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_1798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_21_1840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_21_1874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_1963 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_1980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_1992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_2003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_234 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_262 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_21_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_590 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_594 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_606 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_21_640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_652 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_21_703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_21_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_21_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_21_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_21_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_21_89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1758 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1762 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_178 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1786 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1864 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1868 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_1874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1898 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_1902 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_1912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1963 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_2008 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_214 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_260 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_22_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_282 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_22_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_22_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_22_370 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_402 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_414 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_22_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_22_565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_22_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_22_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_22_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_22_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_22_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_22_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_22_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_22_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_1598 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1678 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1702 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1714 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_2006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_362 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_23_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_402 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_462 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_466 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_23_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_23_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_23_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_73 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_23_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_23_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_23_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_1781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_1928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1948 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_1952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_2005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_2023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_2032 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_2055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_2080 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2095 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_2119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_2243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_2275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_2299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_2304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_2320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_2328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_2335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_2347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_24_264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_24_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_24_717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_24_733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_24_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_24_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_24_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1834 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_1846 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_1907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_1993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2051 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_2066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2070 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_2076 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_2080 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2084 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_2167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_2226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_2230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_2263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_2270 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_2279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_2326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_2335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_408 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_428 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_516 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_520 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_532 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_544 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_25_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_25_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_25_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_25_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_25_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_25_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_25_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_1571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_1780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1792 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_1800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_1856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_1947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_1962 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_1966 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_2027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2046 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_2119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_2251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_2257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_2326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_2334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_2358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_292 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_26_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_568 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_58 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_580 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_639 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_26_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_26_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_26_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_26_726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_730 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_26_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_26_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_13 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1686 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_1738 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1772 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_1852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1868 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_1891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1955 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_2028 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2032 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2052 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2079 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_2088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2092 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_2111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_2167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_2219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_2223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_2299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_2326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_2335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_2359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_25 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_37 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_423 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_49 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_540 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_544 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_27_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_27_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_27_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_27_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_27_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_74 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_27_86 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_27_98 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1052 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_1976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_1980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2196 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_2200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_2301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_2304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_2329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_2341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_486 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_66 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_28_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_834 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_28_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_28_882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_28_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_28_964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_28_968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_28_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1724 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1759 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1879 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_2024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2028 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2040 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2052 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2064 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_2104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_2215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_2232 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_2287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_2312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_2318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_2346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_414 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_568 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_572 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_596 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_638 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_654 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_74 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_746 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_29_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_29_815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_29_830 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_29_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_29_95 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_29_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_29_99 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_10 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1004 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1026 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1074 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1078 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1082 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1214 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1292 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1338 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_134 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1360 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1364 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_138 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_14 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1404 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1504 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1516 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1610 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1622 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1636 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1644 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1678 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1684 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_176 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1762 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1796 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1814 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1858 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1864 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1868 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1888 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_1907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1920 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1970 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1975 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_1984 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_1993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_1996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_20 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_2012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2016 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2020 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2028 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2042 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_2058 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_2079 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_2147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2182 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2232 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2236 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_2244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_2279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_2283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_2299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_2314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_2343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_24 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_338 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_35 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_43 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_452 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_498 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_514 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_578 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_59 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_6 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_626 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_63 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_68 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_730 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_764 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_822 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_830 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_844 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_2_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_2_957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_2_969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_2_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_2_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_2_992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_2_996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1018 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1182 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1254 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_1279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1352 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_1435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_168 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1700 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_2005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_2022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2026 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2038 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_2058 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2074 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2086 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_2117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_2220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_2280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_2284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_316 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_398 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_436 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_30_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_59 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_611 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_622 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_634 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_67 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_786 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_906 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_910 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_922 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_30_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_30_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_30_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_30_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_30_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_30_994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1224 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1700 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1728 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_1740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1772 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1784 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_1881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_204 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_2050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_2070 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_2123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_2173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_2275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_2283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_612 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_63 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_67 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_788 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_792 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_80 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_31_804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_812 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_31_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_31_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_88 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_31_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_31_901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_31_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_31_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1018 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1070 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1082 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1395 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1438 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1462 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1646 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1675 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_1962 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1966 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_1972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_1976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_2027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_2112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_2128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_2300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_414 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_49 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_58 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_684 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_696 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_32_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_32_89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_32_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_32_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_32_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_32_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_32_994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1168 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1370 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1590 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1594 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1598 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1610 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1622 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_1996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_2087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_2108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_2118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2159 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_216 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_2301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_552 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_33_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_712 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_73 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_796 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_33_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_872 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_33_963 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_33_971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_33_978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_33_982 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_33_994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1086 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1158 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1246 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1258 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1286 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1290 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1572 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1576 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_1660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1664 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1832 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1872 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_1912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_1916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_1974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_1977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2078 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_2096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_2219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_2228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_282 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_386 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_398 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_34_62 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_66 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_34_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_738 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_852 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_34_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_34_911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_922 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_34_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_34_987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_34_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1004 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1095 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_1977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_1993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_2032 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2095 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_212 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_2229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_276 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_292 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_340 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_552 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_718 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_764 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_79 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_35_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_87 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_35_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_906 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_35_92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_926 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_35_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_96 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_35_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_35_972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_35_987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1019 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1158 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1186 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1234 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1496 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_1608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1612 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1624 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1636 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1648 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_1672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1700 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_1948 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_1992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_1996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2092 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_2231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_2234 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2246 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2258 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_2266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_2291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_362 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_408 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_463 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_59 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_600 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_616 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_624 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_36_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_80 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_835 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_36_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_36_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_36_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_36_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_36_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_36_995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1002 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_1107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_1206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_1262 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_1524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_1536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_1580 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1596 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1712 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1728 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_1994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_1998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2010 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_2147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_2151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2236 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_2304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_2308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_2344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_438 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_37_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_532 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_540 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_614 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_758 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_37_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_820 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_832 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_37_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_37_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_37_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_37_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_37_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_1010 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1034 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1138 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_1303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1420 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1424 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1732 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1872 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_1930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_2016 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2020 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_2067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_2115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_2217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_2227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_2245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_680 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_687 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_708 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_712 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_724 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_736 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_748 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_38_761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_788 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_792 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_38_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_38_901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_906 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_38_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_38_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_38_986 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_38_998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1031 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1051 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1056 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_1071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_1096 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1668 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1728 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1872 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1888 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_39_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_634 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_638 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_662 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_39_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_39_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_39_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_39_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_39_916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_940 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_39_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1002 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1056 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1282 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1286 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1370 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1382 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1423 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1466 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1506 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_1734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1914 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1926 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_1977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_1980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_1992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2004 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_2008 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_2051 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2070 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_2104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_2160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2182 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_2210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_2234 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_2348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_3_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_374 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_390 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_423 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_45 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_64 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_68 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_80 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_3_815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_3_866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_3_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_3_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_3_972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_984 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_3_996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1078 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_1302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_1328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_40_1376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1404 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1416 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_1517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_40_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_2089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_2150 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_2154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_736 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_752 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_40_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_40_790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_794 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_40_820 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_824 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_848 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_40_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_40_941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_40_954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_970 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_40_978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_40_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_40_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1006 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_41_1239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1356 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1360 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_1489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_1916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1920 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_41_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_2066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2316 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_2320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_2344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_41_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_700 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_708 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_41_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_41_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_41_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_41_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_924 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_41_970 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_41_974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_986 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_41_998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_42_1162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1166 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1178 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1451 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_42_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_1907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_42_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_42_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_42_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_42_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_42_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_42_997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_43_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_43_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_43_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1076 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_43_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_43_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_1293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_43_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_1387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2059 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_2067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_43_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_43_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_43_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_43_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_43_778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_43_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_43_891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_43_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_43_905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_43_912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_43_916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_928 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_940 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_43_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_44_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_44_1114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_44_1124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1176 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_44_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1254 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_44_1280 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_44_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_1454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1466 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1478 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_44_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_44_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_44_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_44_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_44_826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_830 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_842 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_854 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_44_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_44_936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_44_940 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_952 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_44_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_44_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_45_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_1136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_45_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_45_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_2066 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_45_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_45_2320 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_2324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_2328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2340 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_45_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_45_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_45_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_45_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_904 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_45_947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_45_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_45_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_45_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_1108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_1131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_1276 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1300 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_1444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1480 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_46_2285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_46_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_46_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_2329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_46_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_46_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_46_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_46_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_46_933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_46_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_46_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_46_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_46_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_10 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_47_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1084 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_47_1150 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1166 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_1174 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1336 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_22 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2222 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_47_2313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_47_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_34 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_46 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_6 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_47_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_47_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_47_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_47_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_47_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_47_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_48_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_48_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1794 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1818 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_1964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_1980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_48_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_48_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2064 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2076 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_2118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_48_2145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_2149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_2230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2254 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_48_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_50 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_48_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_48_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_66 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_78 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_48_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_48_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_48_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_1094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1554 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_49_1734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_1769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1902 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_1921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_2034 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_2038 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_2089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_2093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_2302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_2327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_2361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_49_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_49_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_49_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_49_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_49_901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_49_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_49_989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1027 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_1042 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_1047 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1079 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1292 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1462 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1535 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_1545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1620 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1716 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1732 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1857 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2068 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2080 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2092 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_2154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_2228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2240 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_2257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_2355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_546 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_56 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_60 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_654 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_694 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_738 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_4_742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_750 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_790 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_4_810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_4_873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_4_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_4_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_4_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_4_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1526 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1678 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1784 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1788 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1818 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_182 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2016 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2020 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_2055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_2063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2095 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_2142 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_2154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_2161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2179 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_50_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_23 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_2310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_2329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_2357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_2360 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_284 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_296 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_354 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_492 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_514 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_518 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_50_528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_50_538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_546 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_574 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_50_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_50_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_50_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_50_993 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1040 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1056 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1184 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1196 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1275 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1302 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1326 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1370 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_1378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_1384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1432 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1436 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1448 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1504 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1508 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1523 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1532 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1544 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1576 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1588 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1611 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_164 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1644 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1648 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1672 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1750 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1760 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1764 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1780 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1784 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1840 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1858 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_188 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_1938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1968 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_198 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1980 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_1991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_1994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_1998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2002 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_2008 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2026 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2030 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_2036 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2040 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2044 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_2050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_2060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_2137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2142 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_2162 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2201 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2216 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_2238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_23 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_2328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_2336 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_2344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_318 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_324 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_358 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_362 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_366 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_37 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_376 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_380 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_386 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_45 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_458 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_478 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_48 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_486 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_52 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_542 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_546 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_594 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_600 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_632 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_644 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_656 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_668 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_71 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_792 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_804 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_51_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_87 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_894 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_51_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_90 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_95 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_51_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_51_966 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_51_978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_986 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_51_992 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_51_995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_52_1000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1011 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1020 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_52_1026 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1058 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1062 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1078 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1082 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1142 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1156 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1171 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1180 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1200 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1214 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1252 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1258 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1272 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1276 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1330 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1334 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1354 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1368 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1388 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1392 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_14 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1407 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1412 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_52_1418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1470 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1494 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1534 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1552 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1572 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1592 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1626 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1630 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1644 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1658 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1662 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1680 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1684 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1722 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1726 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1746 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1782 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1806 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1810 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1814 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1842 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1846 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1862 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1870 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1886 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1891 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1926 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1930 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1946 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_1964 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_1969 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_1978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1984 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_1998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2002 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2042 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2050 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2056 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2060 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2076 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2080 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2094 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2138 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_2167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2191 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2196 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_52_2202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2244 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2254 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2263 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2274 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_2289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_23 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2312 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2316 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_232 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_2322 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2332 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2336 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_2346 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_2350 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_278 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_290 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_33 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_336 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_372 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_38 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_382 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_396 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_400 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_410 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_52_450 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_463 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_468 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_472 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_599 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_604 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_628 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_64 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_666 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_682 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_686 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_690 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_706 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_710 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_715 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_744 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_750 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_764 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_768 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_788 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_802 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_808 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_822 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_826 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_860 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_866 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_880 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_884 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_9 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_91 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_913 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_918 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_932 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_936 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_947 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_96 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_962 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_52_976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_52_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_52_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_52_996 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1016 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1034 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1052 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1146 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1168 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1226 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1248 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1306 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1328 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1342 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1350 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1364 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1386 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1408 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1444 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1519 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1538 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1547 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1575 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1611 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1698 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1720 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1734 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1742 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1756 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1771 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1800 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1818 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1836 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1894 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1911 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1916 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1967 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_1974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_1981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2010 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2032 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2054 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2083 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2134 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2148 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2170 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2228 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_2235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2245 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2308 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_362 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_440 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_458 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_464 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_487 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_493 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_498 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_522 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_551 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_558 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_580 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_602 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_62 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_624 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_638 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_662 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_696 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_718 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_740 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_798 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_834 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_856 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_914 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_950 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_958 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_53_972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_53_987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_53_994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1005 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1154 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1160 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1172 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1192 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1196 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1246 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1256 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1262 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1266 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1270 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1282 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1354 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1474 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1478 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1482 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1486 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1490 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1502 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1510 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1540 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_1563 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1566 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1593 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1605 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1661 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1773 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_181 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1823 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1879 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1882 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1894 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_1902 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_1997 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2071 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2073 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2085 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2097 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2209 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2221 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2239 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_2249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2260 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_2264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2276 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2288 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_2345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_2351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_2359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_381 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_384 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_641 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_754 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_758 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_762 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_770 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_829 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_5_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_5_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_90 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_5_915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_94 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_5_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_5_977 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_5_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_994 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_5_998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1000 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1024 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1048 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1089 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1251 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1340 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1344 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1348 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1352 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1437 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1446 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1521 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1548 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1568 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1572 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1608 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1612 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1616 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1622 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1626 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1630 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1650 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1677 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1703 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1801 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_1837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1885 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1965 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_197 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_1975 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_1979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_2025 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_2043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_206 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2081 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2093 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_2099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_2136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_2140 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2152 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_2175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_2178 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_218 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2202 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_2210 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_2235 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2247 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_2267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_230 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_2323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_2359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_2363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_250 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_289 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_301 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_345 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_409 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_469 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_581 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_637 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_640 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_657 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_681 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_745 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_769 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_781 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_6_896 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_900 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_904 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_6_920 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_941 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_956 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_960 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_6_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_6_972 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_6_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_6_985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_6_988 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_10 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1021 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1033 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1037 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1049 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1065 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1077 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1088 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1145 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1149 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1161 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1189 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_7_1193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1203 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1217 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1233 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1257 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1273 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1294 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1298 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1304 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1310 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1314 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1317 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1329 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1357 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1373 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1385 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1401 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1413 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1426 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1429 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1442 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1446 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1454 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1457 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_1481 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1485 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1497 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1513 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1553 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1562 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1569 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_1577 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1582 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1586 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1590 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1597 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1609 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1618 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1625 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1633 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_165 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1653 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1665 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1674 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_1688 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_1692 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1704 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_7_1709 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1721 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1737 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1749 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1765 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_177 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_1777 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1789 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1793 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1805 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1817 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1821 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1833 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1849 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1861 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1877 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1889 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1905 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1917 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1929 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1933 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_194 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_1945 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_1985 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_1989 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2001 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2013 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2017 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2045 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2057 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_2069 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_207 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2086 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2090 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_2098 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2141 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_2153 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2157 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2169 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_2183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_2185 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_2193 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_22 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_2208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_2213 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_223 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_2241 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2269 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2297 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2325 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_2349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_2353 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_237 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_249 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_281 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_293 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_305 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_309 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_321 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_337 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_349 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_365 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_377 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_393 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_405 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_421 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_433 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_449 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_461 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_477 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_489 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_49 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_501 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_505 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_529 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_533 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_573 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_585 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_589 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_6 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_601 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_617 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_629 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_642 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_645 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_701 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_713 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_73 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_741 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_757 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_772 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_776 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_7_785 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_797 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_813 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_825 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_837 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_841 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_853 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_865 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_869 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_88 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_881 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_897 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_909 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_921 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_7_925 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_937 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_7_949 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_7_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_96 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_970 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_7_981 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_7_999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1015 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1019 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1023 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_1029 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1041 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1053 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1061 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1063 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1075 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1099 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1143 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1155 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1167 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1173 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1205 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1208 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1220 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_8_1225 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_1229 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1243 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1255 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1267 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1285 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1287 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1299 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1311 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1323 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1341 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1367 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1379 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1397 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1430 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1434 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1455 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1467 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1479 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1491 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1509 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_1517 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1525 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1528 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1534 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1537 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1561 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_1565 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1603 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1621 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1647 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1676 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_8_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1689 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1693 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1717 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1729 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_1733 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_1767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_8_1791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1815 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1827 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1845 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1859 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1871 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1883 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1901 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1903 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1915 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1927 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1939 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_1957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_1959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1971 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1983 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_1995 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_265 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_277 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_279 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_291 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_333 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_335 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_347 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_359 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_371 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_389 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_391 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_403 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_415 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_439 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_445 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_459 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_471 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_503 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_515 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_527 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_541 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_545 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_549 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_557 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_559 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_571 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_583 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_613 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_615 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_627 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_8_631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_655 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_659 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_669 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_671 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_683 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_695 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_725 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_727 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_739 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_751 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_774 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_778 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_783 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_795 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_807 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_816 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_820 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_832 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_839 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_8_893 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_895 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_907 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_919 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_931 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_943 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_8_948 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_951 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_959 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_8_962 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_974 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_8_982 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_8_986 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_8_998 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1003 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1009 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1012 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_1022 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1035 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1039 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1043 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1055 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1067 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1079 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_1087 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1091 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_1123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1144 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1147 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1151 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1163 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1175 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1183 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1187 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1190 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1195 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1199 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1211 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1215 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1219 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1227 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1231 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1238 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1242 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1246 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1259 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1313 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1315 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1327 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1339 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1351 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1369 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1378 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1382 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1394 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1406 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1418 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1422 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1425 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1427 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1435 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1443 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1447 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1456 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1460 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1464 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1476 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1483 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1495 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_1499 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1507 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1511 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1516 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1520 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1530 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1536 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1539 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1543 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1555 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1567 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1579 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1591 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_1595 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1607 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1619 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1631 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1649 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1651 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1660 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1664 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1670 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1673 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1685 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_1705 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1707 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1719 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1731 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1743 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1761 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1763 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1775 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1787 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1799 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1808 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1812 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1831 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1867 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1873 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_1875 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1887 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1899 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1908 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1912 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1924 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_1934 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1938 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_1942 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1954 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1966 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1978 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_1987 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_1999 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_2007 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_253 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_261 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_264 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_268 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_271 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_283 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_295 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_303 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_307 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_319 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_331 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_343 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_355 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_361 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_363 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_375 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_383 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_387 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_399 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_411 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_417 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_419 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_431 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_441 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_453 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_465 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_473 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_475 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_484 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_488 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_500 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_512 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_524 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_531 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_535 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_550 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_556 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_560 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_564 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_576 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_584 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_587 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_599 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_611 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_623 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_635 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_638 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_643 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_663 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_667 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_679 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_691 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_697 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_699 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_711 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_723 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_735 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_747 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_753 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_755 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_767 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_779 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_791 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_803 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_6
XFILLER_9_809 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_811 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_819 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_828 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_832 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_4
XFILLER_9_838 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_843 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_847 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_851 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_855 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_863 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XFILLER_9_874 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_878 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_890 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_902 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_914 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_923 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_935 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_8
XFILLER_9_953 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_957 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_961 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_973 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_1
XFILLER_9_976 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__FILL_2
XFILLER_9_979 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XFILLER_9_991 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_12
XPHY_0 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_1 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_10 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_100 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_101 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_102 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_103 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_104 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_105 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_106 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_107 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_108 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_109 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_11 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_110 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_111 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_112 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_113 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_114 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_115 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_116 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_117 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_118 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_119 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_12 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_120 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_121 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_122 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_123 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_124 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_125 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_126 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_127 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_128 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_129 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_13 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_130 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_131 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_132 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_133 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_134 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_135 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_136 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_137 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_138 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_139 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_14 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_15 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_16 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_17 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_18 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_19 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_2 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_20 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_21 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_22 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_23 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_24 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_25 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_26 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_27 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_28 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_29 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_3 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_30 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_31 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_32 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_33 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_34 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_35 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_36 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_37 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_38 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_39 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_4 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_40 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_41 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_42 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_43 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_44 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_45 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_46 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_47 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_48 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_49 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_5 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_50 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_51 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_52 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_53 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_54 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_55 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_56 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_57 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_58 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_59 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_6 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_60 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_61 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_62 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_63 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_64 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_65 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_66 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_67 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_68 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_69 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_7 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_70 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_71 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_72 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_73 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_74 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_75 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_76 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_77 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_78 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_79 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_8 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_80 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_81 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_82 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_83 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_84 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_85 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_86 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_87 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_88 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_89 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_9 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_90 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_91 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_92 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_93 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_94 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_95 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_96 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_97 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_98 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XPHY_99 VSSD VSSD VCCD VCCD SKY130_FD_SC_HD__DECAP_3
XTAP_1000 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1001 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1002 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1003 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1004 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1005 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1006 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1007 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1008 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1009 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1010 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1011 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1012 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1013 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1014 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1015 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1016 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1017 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1018 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1019 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1020 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1021 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1022 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1023 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1024 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1025 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1026 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1027 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1028 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1029 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1030 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1031 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1032 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1033 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1034 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1035 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1036 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1037 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1038 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1039 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1040 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1041 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1042 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1043 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1044 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1045 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1046 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1047 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1048 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1049 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1050 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1051 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1052 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1053 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1054 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1055 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1056 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1057 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1058 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1059 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1060 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1061 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1062 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1063 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1064 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1065 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1066 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1067 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1068 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1069 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1070 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1071 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1072 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1073 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1074 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1075 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1076 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1077 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1078 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1079 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1080 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1081 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1082 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1083 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1084 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1085 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1086 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1087 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1088 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1089 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1090 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1091 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1092 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1093 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1094 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1095 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1096 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1097 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1098 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1099 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1100 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1101 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1102 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1103 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1104 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1105 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1106 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1107 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1108 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1109 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1110 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1111 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1112 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1113 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1114 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1115 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1116 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1117 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1118 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1119 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1120 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1121 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1122 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1123 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1124 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1125 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1126 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1127 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1128 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1129 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1130 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1131 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1132 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1133 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1134 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1135 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1136 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1137 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1138 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1139 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1140 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1141 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1142 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1143 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1144 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1145 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1146 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1147 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1148 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1149 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1150 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1151 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1152 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1153 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1154 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1155 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1156 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1157 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1158 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1159 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1160 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1161 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1162 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1163 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1164 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1165 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1166 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1167 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1168 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1169 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1170 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1171 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1172 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1173 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1174 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1175 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1176 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1177 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1178 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1179 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1180 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1181 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1182 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1183 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1184 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1185 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1186 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1187 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1188 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1189 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1190 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1191 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1192 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1193 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1194 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1195 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1196 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1197 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1198 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1199 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1200 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1201 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1202 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1203 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1204 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1205 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1206 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1207 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1208 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1209 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1210 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1211 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1212 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1213 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1214 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1215 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1216 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1217 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1218 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1219 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1220 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1221 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1222 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1223 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1224 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1225 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1226 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1227 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1228 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1229 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1230 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1231 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1232 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1233 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1234 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1235 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1236 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1237 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1238 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1239 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1240 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1241 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1242 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1243 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1244 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1245 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1246 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1247 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1248 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1249 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1250 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1251 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1252 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1253 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1254 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1255 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1256 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1257 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1258 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1259 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1260 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1261 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1262 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1263 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1264 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1265 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1266 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1267 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1268 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1269 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1270 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1271 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1272 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1273 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1274 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1275 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1276 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1277 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1278 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1279 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1280 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1281 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1282 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1283 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1284 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1285 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1286 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1287 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1288 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1289 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1290 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1291 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1292 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1293 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1294 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1295 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1296 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1297 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1298 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1299 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1300 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1301 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1302 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1303 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1304 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1305 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1306 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1307 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1308 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1309 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1310 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1311 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1312 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1313 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1314 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1315 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1316 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1317 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1318 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1319 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1320 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1321 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1322 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1323 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1324 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1325 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1326 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1327 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1328 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1329 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1330 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1331 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1332 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1333 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1334 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1335 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1336 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1337 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1338 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1339 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1340 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1341 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1342 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1343 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1344 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1345 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1346 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1347 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1348 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1349 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1350 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1351 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1352 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1353 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1354 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1355 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1356 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1357 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1358 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1359 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1360 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1361 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1362 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1363 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1364 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1365 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1366 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1367 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1368 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1369 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1370 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1371 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1372 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1373 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1374 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1375 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1376 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1377 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1378 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1379 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1380 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1381 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1382 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1383 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1384 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1385 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1386 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1387 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1388 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1389 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1390 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1391 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1392 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1393 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1394 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1395 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1396 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1397 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1398 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1399 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_140 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1400 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1401 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1402 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1403 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1404 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1405 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1406 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1407 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1408 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1409 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_141 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1410 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1411 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1412 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1413 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1414 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1415 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1416 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1417 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1418 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1419 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_142 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1420 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1421 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1422 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1423 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1424 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1425 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1426 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1427 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1428 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1429 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_143 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1430 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1431 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1432 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1433 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1434 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1435 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1436 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1437 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1438 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1439 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_144 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1440 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1441 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1442 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1443 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1444 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1445 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1446 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1447 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1448 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1449 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_145 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1450 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1451 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1452 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1453 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1454 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1455 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1456 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1457 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1458 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1459 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_146 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1460 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1461 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1462 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1463 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1464 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1465 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1466 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1467 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1468 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1469 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_147 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1470 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1471 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1472 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1473 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1474 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1475 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1476 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1477 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1478 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1479 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_148 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1480 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1481 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1482 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1483 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1484 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1485 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1486 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1487 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1488 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1489 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_149 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1490 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1491 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1492 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1493 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1494 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1495 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1496 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1497 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1498 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1499 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_150 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1500 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1501 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1502 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1503 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1504 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1505 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1506 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1507 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1508 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1509 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_151 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1510 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1511 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1512 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1513 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1514 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1515 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1516 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1517 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1518 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1519 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_152 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1520 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1521 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1522 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1523 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1524 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1525 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1526 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1527 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1528 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1529 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_153 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1530 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1531 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1532 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1533 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1534 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1535 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1536 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1537 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1538 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1539 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_154 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1540 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1541 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1542 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1543 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1544 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1545 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1546 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1547 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1548 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1549 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_155 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1550 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1551 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1552 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1553 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1554 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1555 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1556 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1557 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1558 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1559 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_156 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1560 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1561 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1562 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1563 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1564 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1565 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1566 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1567 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1568 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1569 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_157 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1570 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1571 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1572 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1573 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1574 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1575 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1576 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1577 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1578 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1579 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_158 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1580 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1581 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1582 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1583 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1584 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1585 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1586 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1587 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1588 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1589 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_159 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1590 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1591 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1592 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1593 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1594 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1595 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1596 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1597 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1598 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1599 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_160 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1600 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1601 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1602 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1603 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1604 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1605 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1606 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1607 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1608 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1609 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_161 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1610 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1611 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1612 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1613 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1614 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1615 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1616 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1617 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1618 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1619 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_162 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1620 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1621 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1622 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1623 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1624 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1625 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1626 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1627 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1628 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1629 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_163 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1630 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1631 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1632 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1633 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1634 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1635 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1636 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1637 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1638 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1639 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_164 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1640 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1641 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1642 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1643 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1644 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1645 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1646 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1647 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1648 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1649 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_165 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1650 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1651 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1652 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1653 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1654 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1655 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1656 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1657 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1658 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1659 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_166 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1660 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1661 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1662 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1663 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1664 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1665 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1666 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1667 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1668 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1669 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_167 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1670 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1671 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1672 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1673 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1674 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1675 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1676 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1677 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1678 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1679 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_168 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1680 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1681 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1682 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1683 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1684 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1685 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1686 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1687 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1688 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1689 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_169 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1690 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1691 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1692 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1693 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1694 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1695 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1696 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1697 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1698 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1699 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_170 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1700 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1701 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1702 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1703 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1704 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1705 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1706 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1707 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1708 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1709 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_171 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1710 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1711 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1712 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1713 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1714 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1715 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1716 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1717 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1718 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1719 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_172 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1720 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1721 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1722 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1723 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1724 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1725 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1726 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1727 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1728 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1729 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_173 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1730 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1731 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1732 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1733 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1734 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1735 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1736 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1737 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1738 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1739 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_174 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1740 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1741 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1742 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1743 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1744 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1745 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1746 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1747 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1748 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1749 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_175 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1750 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1751 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1752 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1753 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1754 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1755 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1756 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1757 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1758 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1759 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_176 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1760 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1761 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1762 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1763 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1764 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1765 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1766 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1767 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1768 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1769 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_177 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1770 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1771 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1772 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1773 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1774 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1775 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1776 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1777 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1778 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1779 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_178 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1780 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1781 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1782 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1783 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1784 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1785 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1786 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1787 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1788 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1789 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_179 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1790 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1791 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1792 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1793 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1794 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1795 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1796 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1797 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1798 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1799 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_180 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1800 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1801 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1802 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1803 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1804 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1805 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1806 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1807 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1808 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1809 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_181 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1810 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1811 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1812 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1813 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1814 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1815 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1816 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1817 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1818 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1819 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_182 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1820 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1821 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1822 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1823 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1824 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1825 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1826 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1827 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1828 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1829 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_183 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1830 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1831 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1832 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1833 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1834 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1835 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1836 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1837 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1838 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1839 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_184 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1840 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1841 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1842 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1843 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1844 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1845 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1846 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1847 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1848 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1849 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_185 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1850 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1851 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1852 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1853 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1854 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1855 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1856 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1857 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1858 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1859 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_186 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1860 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1861 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1862 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1863 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1864 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1865 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1866 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1867 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1868 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1869 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_187 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1870 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1871 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1872 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1873 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1874 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1875 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1876 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1877 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1878 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1879 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_188 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1880 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1881 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1882 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1883 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1884 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1885 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1886 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1887 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1888 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1889 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_189 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1890 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1891 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1892 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1893 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1894 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1895 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1896 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1897 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1898 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1899 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_190 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1900 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1901 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1902 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1903 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1904 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1905 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1906 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1907 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1908 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1909 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_191 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1910 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1911 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1912 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1913 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1914 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1915 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1916 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1917 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1918 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1919 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_192 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1920 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1921 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1922 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1923 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1924 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1925 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1926 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1927 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1928 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1929 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_193 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1930 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1931 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1932 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1933 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1934 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1935 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1936 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1937 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1938 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1939 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_194 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1940 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1941 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1942 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1943 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1944 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1945 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1946 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1947 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1948 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1949 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_195 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1950 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1951 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1952 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1953 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1954 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1955 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1956 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1957 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1958 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1959 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_196 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1960 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1961 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1962 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1963 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1964 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1965 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1966 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1967 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1968 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1969 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_197 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1970 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1971 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1972 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1973 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1974 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1975 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1976 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1977 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1978 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1979 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_198 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1980 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1981 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1982 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1983 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1984 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1985 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1986 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1987 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1988 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1989 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_199 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1990 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1991 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1992 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1993 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1994 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1995 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1996 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1997 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1998 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_1999 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_200 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2000 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2001 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2002 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2003 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2004 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2005 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2006 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2007 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2008 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2009 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_201 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2010 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2011 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2012 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2013 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2014 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2015 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2016 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2017 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2018 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2019 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_202 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2020 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2021 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2022 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2023 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2024 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2025 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2026 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2027 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2028 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2029 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_203 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2030 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2031 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2032 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2033 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2034 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2035 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2036 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2037 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2038 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2039 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_204 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2040 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2041 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2042 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2043 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2044 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2045 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2046 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2047 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2048 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2049 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_205 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2050 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2051 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2052 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2053 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2054 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2055 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2056 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2057 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2058 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2059 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_206 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2060 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2061 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2062 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2063 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2064 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2065 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2066 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2067 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2068 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2069 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_207 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2070 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2071 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2072 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2073 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2074 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2075 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2076 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2077 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2078 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2079 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_208 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2080 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2081 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2082 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2083 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2084 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2085 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2086 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2087 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2088 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2089 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_209 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2090 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2091 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2092 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2093 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2094 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2095 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2096 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2097 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2098 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2099 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_210 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2100 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2101 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2102 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2103 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2104 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2105 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2106 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2107 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2108 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2109 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_211 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2110 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2111 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2112 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2113 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2114 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2115 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2116 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2117 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2118 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2119 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_212 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2120 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2121 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2122 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2123 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2124 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2125 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2126 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2127 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2128 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2129 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_213 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2130 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2131 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2132 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2133 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2134 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2135 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2136 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2137 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2138 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2139 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_214 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2140 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2141 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2142 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2143 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2144 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2145 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2146 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2147 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2148 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2149 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_215 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2150 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2151 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2152 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2153 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2154 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2155 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2156 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2157 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2158 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2159 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_216 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2160 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2161 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2162 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2163 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2164 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2165 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2166 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2167 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2168 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2169 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_217 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2170 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2171 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2172 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2173 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2174 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2175 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2176 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2177 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2178 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2179 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_218 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2180 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2181 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2182 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2183 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2184 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2185 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2186 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2187 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2188 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2189 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_219 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2190 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2191 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2192 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2193 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2194 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2195 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2196 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2197 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2198 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2199 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_220 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2200 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2201 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2202 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2203 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2204 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2205 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2206 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2207 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2208 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2209 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_221 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2210 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2211 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2212 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2213 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2214 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2215 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2216 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2217 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2218 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2219 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_222 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2220 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2221 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2222 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2223 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2224 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2225 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2226 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2227 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2228 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2229 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_223 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2230 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2231 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2232 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2233 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2234 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2235 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2236 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2237 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2238 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2239 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_224 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2240 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2241 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2242 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2243 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2244 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2245 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2246 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2247 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2248 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2249 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_225 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2250 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2251 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2252 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2253 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2254 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2255 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2256 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2257 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2258 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2259 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_226 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2260 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2261 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2262 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2263 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2264 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2265 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2266 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2267 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2268 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_2269 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_227 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_228 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_229 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_230 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_231 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_232 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_233 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_234 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_235 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_236 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_237 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_238 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_239 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_240 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_241 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_242 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_243 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_244 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_245 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_246 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_247 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_248 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_249 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_250 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_251 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_252 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_253 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_254 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_255 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_256 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_257 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_258 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_259 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_260 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_261 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_262 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_263 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_264 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_265 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_266 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_267 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_268 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_269 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_270 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_271 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_272 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_273 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_274 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_275 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_276 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_277 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_278 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_279 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_280 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_281 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_282 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_283 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_284 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_285 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_286 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_287 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_288 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_289 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_290 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_291 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_292 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_293 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_294 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_295 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_296 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_297 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_298 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_299 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_300 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_301 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_302 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_303 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_304 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_305 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_306 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_307 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_308 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_309 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_310 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_311 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_312 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_313 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_314 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_315 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_316 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_317 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_318 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_319 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_320 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_321 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_322 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_323 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_324 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_325 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_326 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_327 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_328 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_329 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_330 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_331 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_332 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_333 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_334 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_335 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_336 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_337 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_338 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_339 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_340 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_341 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_342 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_343 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_344 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_345 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_346 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_347 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_348 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_349 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_350 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_351 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_352 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_353 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_354 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_355 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_356 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_357 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_358 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_359 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_360 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_361 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_362 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_363 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_364 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_365 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_366 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_367 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_368 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_369 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_370 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_371 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_372 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_373 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_374 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_375 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_376 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_377 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_378 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_379 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_380 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_381 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_382 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_383 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_384 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_385 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_386 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_387 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_388 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_389 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_390 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_391 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_392 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_393 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_394 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_395 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_396 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_397 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_398 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_399 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_400 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_401 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_402 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_403 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_404 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_405 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_406 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_407 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_408 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_409 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_410 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_411 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_412 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_413 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_414 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_415 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_416 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_417 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_418 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_419 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_420 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_421 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_422 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_423 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_424 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_425 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_426 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_427 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_428 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_429 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_430 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_431 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_432 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_433 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_434 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_435 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_436 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_437 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_438 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_439 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_440 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_441 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_442 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_443 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_444 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_445 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_446 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_447 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_448 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_449 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_450 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_451 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_452 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_453 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_454 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_455 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_456 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_457 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_458 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_459 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_460 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_461 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_462 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_463 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_464 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_465 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_466 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_467 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_468 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_469 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_470 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_471 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_472 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_473 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_474 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_475 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_476 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_477 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_478 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_479 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_480 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_481 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_482 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_483 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_484 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_485 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_486 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_487 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_488 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_489 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_490 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_491 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_492 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_493 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_494 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_495 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_496 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_497 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_498 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_499 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_500 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_501 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_502 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_503 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_504 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_505 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_506 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_507 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_508 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_509 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_510 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_511 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_512 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_513 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_514 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_515 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_516 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_517 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_518 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_519 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_520 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_521 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_522 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_523 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_524 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_525 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_526 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_527 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_528 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_529 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_530 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_531 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_532 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_533 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_534 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_535 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_536 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_537 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_538 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_539 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_540 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_541 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_542 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_543 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_544 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_545 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_546 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_547 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_548 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_549 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_550 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_551 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_552 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_553 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_554 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_555 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_556 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_557 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_558 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_559 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_560 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_561 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_562 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_563 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_564 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_565 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_566 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_567 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_568 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_569 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_570 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_571 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_572 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_573 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_574 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_575 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_576 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_577 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_578 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_579 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_580 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_581 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_582 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_583 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_584 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_585 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_586 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_587 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_588 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_589 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_590 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_591 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_592 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_593 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_594 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_595 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_596 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_597 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_598 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_599 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_600 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_601 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_602 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_603 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_604 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_605 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_606 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_607 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_608 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_609 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_610 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_611 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_612 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_613 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_614 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_615 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_616 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_617 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_618 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_619 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_620 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_621 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_622 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_623 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_624 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_625 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_626 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_627 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_628 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_629 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_630 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_631 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_632 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_633 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_634 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_635 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_636 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_637 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_638 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_639 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_640 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_641 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_642 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_643 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_644 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_645 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_646 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_647 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_648 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_649 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_650 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_651 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_652 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_653 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_654 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_655 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_656 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_657 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_658 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_659 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_660 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_661 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_662 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_663 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_664 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_665 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_666 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_667 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_668 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_669 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_670 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_671 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_672 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_673 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_674 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_675 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_676 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_677 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_678 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_679 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_680 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_681 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_682 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_683 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_684 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_685 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_686 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_687 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_688 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_689 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_690 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_691 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_692 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_693 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_694 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_695 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_696 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_697 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_698 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_699 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_700 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_701 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_702 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_703 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_704 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_705 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_706 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_707 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_708 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_709 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_710 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_711 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_712 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_713 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_714 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_715 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_716 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_717 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_718 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_719 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_720 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_721 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_722 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_723 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_724 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_725 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_726 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_727 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_728 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_729 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_730 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_731 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_732 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_733 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_734 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_735 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_736 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_737 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_738 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_739 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_740 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_741 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_742 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_743 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_744 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_745 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_746 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_747 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_748 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_749 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_750 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_751 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_752 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_753 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_754 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_755 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_756 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_757 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_758 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_759 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_760 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_761 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_762 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_763 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_764 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_765 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_766 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_767 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_768 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_769 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_770 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_771 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_772 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_773 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_774 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_775 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_776 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_777 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_778 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_779 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_780 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_781 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_782 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_783 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_784 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_785 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_786 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_787 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_788 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_789 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_790 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_791 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_792 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_793 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_794 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_795 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_796 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_797 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_798 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_799 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_800 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_801 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_802 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_803 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_804 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_805 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_806 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_807 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_808 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_809 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_810 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_811 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_812 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_813 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_814 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_815 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_816 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_817 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_818 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_819 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_820 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_821 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_822 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_823 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_824 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_825 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_826 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_827 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_828 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_829 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_830 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_831 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_832 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_833 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_834 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_835 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_836 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_837 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_838 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_839 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_840 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_841 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_842 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_843 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_844 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_845 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_846 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_847 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_848 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_849 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_850 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_851 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_852 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_853 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_854 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_855 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_856 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_857 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_858 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_859 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_860 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_861 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_862 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_863 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_864 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_865 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_866 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_867 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_868 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_869 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_870 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_871 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_872 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_873 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_874 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_875 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_876 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_877 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_878 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_879 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_880 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_881 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_882 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_883 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_884 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_885 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_886 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_887 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_888 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_889 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_890 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_891 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_892 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_893 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_894 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_895 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_896 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_897 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_898 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_899 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_900 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_901 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_902 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_903 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_904 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_905 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_906 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_907 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_908 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_909 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_910 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_911 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_912 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_913 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_914 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_915 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_916 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_917 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_918 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_919 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_920 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_921 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_922 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_923 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_924 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_925 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_926 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_927 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_928 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_929 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_930 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_931 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_932 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_933 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_934 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_935 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_936 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_937 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_938 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_939 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_940 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_941 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_942 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_943 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_944 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_945 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_946 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_947 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_948 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_949 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_950 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_951 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_952 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_953 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_954 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_955 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_956 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_957 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_958 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_959 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_960 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_961 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_962 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_963 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_964 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_965 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_966 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_967 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_968 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_969 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_970 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_971 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_972 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_973 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_974 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_975 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_976 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_977 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_978 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_979 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_980 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_981 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_982 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_983 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_984 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_985 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_986 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_987 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_988 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_989 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_990 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_991 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_992 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_993 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_994 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_995 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_996 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_997 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_998 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_999 VSSD VCCD SKY130_FD_SC_HD__TAPVPWRVGND_1
X_329_ NET478 VSSD VSSD VCCD VCCD _291_ SKY130_FD_SC_HD__INV_2
X_330_ NET479 VSSD VSSD VCCD VCCD _292_ SKY130_FD_SC_HD__CLKINV_2
X_331_ NET480 VSSD VSSD VCCD VCCD _293_ SKY130_FD_SC_HD__CLKINV_2
X_332_ NET481 VSSD VSSD VCCD VCCD _294_ SKY130_FD_SC_HD__CLKINV_2
X_333_ NET483 VSSD VSSD VCCD VCCD _296_ SKY130_FD_SC_HD__INV_2
X_334_ NET484 VSSD VSSD VCCD VCCD _297_ SKY130_FD_SC_HD__INV_2
X_335_ NET485 VSSD VSSD VCCD VCCD _298_ SKY130_FD_SC_HD__INV_2
X_336_ NET486 VSSD VSSD VCCD VCCD _299_ SKY130_FD_SC_HD__INV_2
X_337_ NET487 VSSD VSSD VCCD VCCD _300_ SKY130_FD_SC_HD__INV_2
X_338_ NET488 VSSD VSSD VCCD VCCD _301_ SKY130_FD_SC_HD__INV_2
X_339_ NET489 VSSD VSSD VCCD VCCD _302_ SKY130_FD_SC_HD__INV_2
X_340_ NET490 VSSD VSSD VCCD VCCD _303_ SKY130_FD_SC_HD__INV_2
X_341_ NET491 VSSD VSSD VCCD VCCD _304_ SKY130_FD_SC_HD__INV_2
X_342_ NET492 VSSD VSSD VCCD VCCD _305_ SKY130_FD_SC_HD__INV_2
X_343_ NET494 VSSD VSSD VCCD VCCD _307_ SKY130_FD_SC_HD__INV_2
X_344_ NET495 VSSD VSSD VCCD VCCD _308_ SKY130_FD_SC_HD__INV_2
X_345_ NET496 VSSD VSSD VCCD VCCD _309_ SKY130_FD_SC_HD__INV_2
X_346_ NET497 VSSD VSSD VCCD VCCD _310_ SKY130_FD_SC_HD__INV_2
X_347_ NET498 VSSD VSSD VCCD VCCD _311_ SKY130_FD_SC_HD__INV_2
X_348_ NET499 VSSD VSSD VCCD VCCD _312_ SKY130_FD_SC_HD__INV_2
X_349_ NET500 VSSD VSSD VCCD VCCD _313_ SKY130_FD_SC_HD__INV_2
X_350_ NET501 VSSD VSSD VCCD VCCD _314_ SKY130_FD_SC_HD__INV_2
X_351_ NET502 VSSD VSSD VCCD VCCD _315_ SKY130_FD_SC_HD__INV_2
X_352_ NET503 VSSD VSSD VCCD VCCD _316_ SKY130_FD_SC_HD__INV_2
X_353_ NET505 VSSD VSSD VCCD VCCD _318_ SKY130_FD_SC_HD__INV_2
X_354_ NET506 VSSD VSSD VCCD VCCD _319_ SKY130_FD_SC_HD__INV_2
X_355_ NET507 VSSD VSSD VCCD VCCD _320_ SKY130_FD_SC_HD__INV_2
X_356_ NET508 VSSD VSSD VCCD VCCD _321_ SKY130_FD_SC_HD__INV_2
X_357_ NET509 VSSD VSSD VCCD VCCD _322_ SKY130_FD_SC_HD__INV_2
X_358_ NET510 VSSD VSSD VCCD VCCD _323_ SKY130_FD_SC_HD__INV_2
X_359_ NET511 VSSD VSSD VCCD VCCD _324_ SKY130_FD_SC_HD__INV_2
X_360_ NET512 VSSD VSSD VCCD VCCD _325_ SKY130_FD_SC_HD__INV_2
X_361_ NET513 VSSD VSSD VCCD VCCD _326_ SKY130_FD_SC_HD__INV_2
X_362_ NET514 VSSD VSSD VCCD VCCD _327_ SKY130_FD_SC_HD__CLKINV_2
X_363_ NET389 VSSD VSSD VCCD VCCD _202_ SKY130_FD_SC_HD__INV_2
X_364_ NET390 VSSD VSSD VCCD VCCD _203_ SKY130_FD_SC_HD__INV_2
X_365_ NET391 VSSD VSSD VCCD VCCD _204_ SKY130_FD_SC_HD__INV_2
X_366_ NET392 VSSD VSSD VCCD VCCD _205_ SKY130_FD_SC_HD__INV_2
X_367_ NET393 VSSD VSSD VCCD VCCD _206_ SKY130_FD_SC_HD__INV_2
X_368_ NET394 VSSD VSSD VCCD VCCD _207_ SKY130_FD_SC_HD__INV_2
X_369_ NET395 VSSD VSSD VCCD VCCD _208_ SKY130_FD_SC_HD__INV_2
X_370_ NET396 VSSD VSSD VCCD VCCD _209_ SKY130_FD_SC_HD__INV_2
X_371_ NET397 VSSD VSSD VCCD VCCD _210_ SKY130_FD_SC_HD__INV_2
X_372_ NET398 VSSD VSSD VCCD VCCD _211_ SKY130_FD_SC_HD__INV_2
X_373_ NET400 VSSD VSSD VCCD VCCD _213_ SKY130_FD_SC_HD__INV_2
X_374_ NET401 VSSD VSSD VCCD VCCD _214_ SKY130_FD_SC_HD__INV_2
X_375_ NET402 VSSD VSSD VCCD VCCD _215_ SKY130_FD_SC_HD__INV_2
X_376_ NET403 VSSD VSSD VCCD VCCD _216_ SKY130_FD_SC_HD__INV_2
X_377_ NET404 VSSD VSSD VCCD VCCD _217_ SKY130_FD_SC_HD__INV_2
X_378_ NET405 VSSD VSSD VCCD VCCD _218_ SKY130_FD_SC_HD__INV_2
X_379_ NET406 VSSD VSSD VCCD VCCD _219_ SKY130_FD_SC_HD__INV_2
X_380_ NET407 VSSD VSSD VCCD VCCD _220_ SKY130_FD_SC_HD__INV_2
X_381_ NET408 VSSD VSSD VCCD VCCD _221_ SKY130_FD_SC_HD__INV_2
X_382_ NET409 VSSD VSSD VCCD VCCD _222_ SKY130_FD_SC_HD__INV_2
X_383_ NET411 VSSD VSSD VCCD VCCD _224_ SKY130_FD_SC_HD__INV_2
X_384_ NET412 VSSD VSSD VCCD VCCD _225_ SKY130_FD_SC_HD__INV_2
X_385_ NET413 VSSD VSSD VCCD VCCD _226_ SKY130_FD_SC_HD__INV_2
X_386_ NET414 VSSD VSSD VCCD VCCD _227_ SKY130_FD_SC_HD__INV_2
X_387_ NET415 VSSD VSSD VCCD VCCD _228_ SKY130_FD_SC_HD__INV_2
X_388_ NET416 VSSD VSSD VCCD VCCD _229_ SKY130_FD_SC_HD__INV_2
X_389_ NET417 VSSD VSSD VCCD VCCD _230_ SKY130_FD_SC_HD__INV_2
X_390_ NET418 VSSD VSSD VCCD VCCD _231_ SKY130_FD_SC_HD__INV_2
X_391_ NET1 VSSD VSSD VCCD VCCD _000_ SKY130_FD_SC_HD__INV_2
X_392_ NET2 VSSD VSSD VCCD VCCD _001_ SKY130_FD_SC_HD__INV_4
X_393_ NET549 VSSD VSSD VCCD VCCD _002_ SKY130_FD_SC_HD__INV_6
X_394_ NET619 VSSD VSSD VCCD VCCD _003_ SKY130_FD_SC_HD__CLKINV_4
X_395_ NET620 VSSD VSSD VCCD VCCD _004_ SKY130_FD_SC_HD__CLKINV_2
X_396_ NET615 VSSD VSSD VCCD VCCD _005_ SKY130_FD_SC_HD__INV_2
X_397_ NET616 VSSD VSSD VCCD VCCD _006_ SKY130_FD_SC_HD__INV_2
X_398_ NET617 VSSD VSSD VCCD VCCD _007_ SKY130_FD_SC_HD__INV_2
X_399_ NET618 VSSD VSSD VCCD VCCD _008_ SKY130_FD_SC_HD__INV_2
X_400_ NET517 VSSD VSSD VCCD VCCD _009_ SKY130_FD_SC_HD__INV_2
X_401_ NET528 VSSD VSSD VCCD VCCD _020_ SKY130_FD_SC_HD__INV_12
X_402_ NET539 VSSD VSSD VCCD VCCD _031_ SKY130_FD_SC_HD__INV_2
X_403_ NET542 VSSD VSSD VCCD VCCD _034_ SKY130_FD_SC_HD__INV_12
X_404_ NET543 VSSD VSSD VCCD VCCD _035_ SKY130_FD_SC_HD__INV_2
X_405_ NET544 VSSD VSSD VCCD VCCD _036_ SKY130_FD_SC_HD__INV_12
X_406_ NET545 VSSD VSSD VCCD VCCD _037_ SKY130_FD_SC_HD__CLKINV_8
X_407_ NET546 VSSD VSSD VCCD VCCD _038_ SKY130_FD_SC_HD__INV_12
X_408_ NET547 VSSD VSSD VCCD VCCD _039_ SKY130_FD_SC_HD__INV_12
X_409_ NET548 VSSD VSSD VCCD VCCD _040_ SKY130_FD_SC_HD__INV_6
X_410_ NET518 VSSD VSSD VCCD VCCD _010_ SKY130_FD_SC_HD__CLKINV_2
X_411_ NET519 VSSD VSSD VCCD VCCD _011_ SKY130_FD_SC_HD__INV_6
X_412_ NET520 VSSD VSSD VCCD VCCD _012_ SKY130_FD_SC_HD__INV_8
X_413_ NET521 VSSD VSSD VCCD VCCD _013_ SKY130_FD_SC_HD__INV_6
X_414_ NET522 VSSD VSSD VCCD VCCD _014_ SKY130_FD_SC_HD__CLKINV_8
X_415_ NET523 VSSD VSSD VCCD VCCD _015_ SKY130_FD_SC_HD__INV_12
X_416_ NET524 VSSD VSSD VCCD VCCD _016_ SKY130_FD_SC_HD__INV_12
X_417_ NET525 VSSD VSSD VCCD VCCD _017_ SKY130_FD_SC_HD__INV_6
X_418_ NET526 VSSD VSSD VCCD VCCD _018_ SKY130_FD_SC_HD__INV_12
X_419_ NET527 VSSD VSSD VCCD VCCD _019_ SKY130_FD_SC_HD__INV_8
X_420_ NET529 VSSD VSSD VCCD VCCD _021_ SKY130_FD_SC_HD__CLKINV_8
X_421_ NET530 VSSD VSSD VCCD VCCD _022_ SKY130_FD_SC_HD__INV_12
X_422_ NET531 VSSD VSSD VCCD VCCD _023_ SKY130_FD_SC_HD__CLKINV_8
X_423_ NET532 VSSD VSSD VCCD VCCD _024_ SKY130_FD_SC_HD__INV_8
X_424_ NET533 VSSD VSSD VCCD VCCD _025_ SKY130_FD_SC_HD__INV_12
X_425_ NET534 VSSD VSSD VCCD VCCD _026_ SKY130_FD_SC_HD__CLKINV_8
X_426_ NET535 VSSD VSSD VCCD VCCD _027_ SKY130_FD_SC_HD__INV_8
X_427_ NET536 VSSD VSSD VCCD VCCD _028_ SKY130_FD_SC_HD__INV_8
X_428_ NET537 VSSD VSSD VCCD VCCD _029_ SKY130_FD_SC_HD__INV_8
X_429_ NET538 VSSD VSSD VCCD VCCD _030_ SKY130_FD_SC_HD__CLKINV_8
X_430_ NET540 VSSD VSSD VCCD VCCD _032_ SKY130_FD_SC_HD__CLKINV_8
X_431_ NET541 VSSD VSSD VCCD VCCD _033_ SKY130_FD_SC_HD__CLKINV_8
X_432_ NET582 VSSD VSSD VCCD VCCD _041_ SKY130_FD_SC_HD__INV_6
X_433_ NET593 VSSD VSSD VCCD VCCD _052_ SKY130_FD_SC_HD__INV_4
X_434_ NET604 VSSD VSSD VCCD VCCD _063_ SKY130_FD_SC_HD__CLKINV_4
X_435_ NET607 VSSD VSSD VCCD VCCD _066_ SKY130_FD_SC_HD__INV_4
X_436_ NET608 VSSD VSSD VCCD VCCD _067_ SKY130_FD_SC_HD__INV_4
X_437_ NET609 VSSD VSSD VCCD VCCD _068_ SKY130_FD_SC_HD__INV_4
X_438_ NET610 VSSD VSSD VCCD VCCD _069_ SKY130_FD_SC_HD__INV_4
X_439_ NET611 VSSD VSSD VCCD VCCD _070_ SKY130_FD_SC_HD__INV_4
X_440_ NET612 VSSD VSSD VCCD VCCD _071_ SKY130_FD_SC_HD__CLKINV_4
X_441_ NET613 VSSD VSSD VCCD VCCD _072_ SKY130_FD_SC_HD__INV_6
X_442_ NET583 VSSD VSSD VCCD VCCD _042_ SKY130_FD_SC_HD__INV_4
X_443_ NET584 VSSD VSSD VCCD VCCD _043_ SKY130_FD_SC_HD__CLKINV_4
X_444_ NET585 VSSD VSSD VCCD VCCD _044_ SKY130_FD_SC_HD__INV_4
X_445_ NET586 VSSD VSSD VCCD VCCD _045_ SKY130_FD_SC_HD__INV_2
X_446_ NET587 VSSD VSSD VCCD VCCD _046_ SKY130_FD_SC_HD__INV_2
X_447_ NET588 VSSD VSSD VCCD VCCD _047_ SKY130_FD_SC_HD__INV_4
X_448_ NET589 VSSD VSSD VCCD VCCD _048_ SKY130_FD_SC_HD__INV_6
X_449_ NET590 VSSD VSSD VCCD VCCD _049_ SKY130_FD_SC_HD__CLKINV_4
X_450_ NET591 VSSD VSSD VCCD VCCD _050_ SKY130_FD_SC_HD__INV_6
X_451_ NET592 VSSD VSSD VCCD VCCD _051_ SKY130_FD_SC_HD__INV_6
X_452_ NET594 VSSD VSSD VCCD VCCD _053_ SKY130_FD_SC_HD__INV_4
X_453_ NET595 VSSD VSSD VCCD VCCD _054_ SKY130_FD_SC_HD__INV_6
X_454_ NET596 VSSD VSSD VCCD VCCD _055_ SKY130_FD_SC_HD__INV_4
X_455_ NET597 VSSD VSSD VCCD VCCD _056_ SKY130_FD_SC_HD__INV_4
X_456_ NET598 VSSD VSSD VCCD VCCD _057_ SKY130_FD_SC_HD__INV_6
X_457_ NET599 VSSD VSSD VCCD VCCD _058_ SKY130_FD_SC_HD__INV_4
X_458_ NET600 VSSD VSSD VCCD VCCD _059_ SKY130_FD_SC_HD__INV_6
X_459_ NET601 VSSD VSSD VCCD VCCD _060_ SKY130_FD_SC_HD__CLKINV_4
X_460_ NET602 VSSD VSSD VCCD VCCD _061_ SKY130_FD_SC_HD__INV_4
X_461_ NET603 VSSD VSSD VCCD VCCD _062_ SKY130_FD_SC_HD__INV_4
X_462_ NET605 VSSD VSSD VCCD VCCD _064_ SKY130_FD_SC_HD__INV_4
X_463_ NET606 VSSD VSSD VCCD VCCD _065_ SKY130_FD_SC_HD__CLKINV_4
X_464_ NET132 VSSD VSSD VCCD VCCD _073_ SKY130_FD_SC_HD__CLKINV_2
X_465_ NET171 VSSD VSSD VCCD VCCD _112_ SKY130_FD_SC_HD__INV_2
X_466_ NET182 VSSD VSSD VCCD VCCD _123_ SKY130_FD_SC_HD__CLKINV_2
X_467_ NET193 VSSD VSSD VCCD VCCD _134_ SKY130_FD_SC_HD__CLKINV_2
X_468_ NET204 VSSD VSSD VCCD VCCD _145_ SKY130_FD_SC_HD__CLKINV_2
X_469_ NET215 VSSD VSSD VCCD VCCD _156_ SKY130_FD_SC_HD__INV_2
X_470_ NET226 VSSD VSSD VCCD VCCD _167_ SKY130_FD_SC_HD__CLKINV_2
X_471_ NET237 VSSD VSSD VCCD VCCD _178_ SKY130_FD_SC_HD__CLKINV_2
X_472_ NET248 VSSD VSSD VCCD VCCD _189_ SKY130_FD_SC_HD__CLKINV_2
X_473_ NET259 VSSD VSSD VCCD VCCD _200_ SKY130_FD_SC_HD__INV_2
X_474_ NET143 VSSD VSSD VCCD VCCD _084_ SKY130_FD_SC_HD__INV_2
X_475_ NET154 VSSD VSSD VCCD VCCD _095_ SKY130_FD_SC_HD__CLKINV_2
X_476_ NET163 VSSD VSSD VCCD VCCD _104_ SKY130_FD_SC_HD__CLKINV_2
X_477_ NET164 VSSD VSSD VCCD VCCD _105_ SKY130_FD_SC_HD__INV_2
X_478_ NET165 VSSD VSSD VCCD VCCD _106_ SKY130_FD_SC_HD__INV_2
X_479_ NET166 VSSD VSSD VCCD VCCD _107_ SKY130_FD_SC_HD__CLKINV_2
X_480_ NET167 VSSD VSSD VCCD VCCD _108_ SKY130_FD_SC_HD__CLKINV_2
X_481_ NET168 VSSD VSSD VCCD VCCD _109_ SKY130_FD_SC_HD__INV_2
X_482_ NET169 VSSD VSSD VCCD VCCD _110_ SKY130_FD_SC_HD__INV_2
X_483_ NET170 VSSD VSSD VCCD VCCD _111_ SKY130_FD_SC_HD__INV_2
X_484_ NET172 VSSD VSSD VCCD VCCD _113_ SKY130_FD_SC_HD__INV_2
X_485_ NET173 VSSD VSSD VCCD VCCD _114_ SKY130_FD_SC_HD__INV_2
X_486_ NET174 VSSD VSSD VCCD VCCD _115_ SKY130_FD_SC_HD__CLKINV_2
X_487_ NET175 VSSD VSSD VCCD VCCD _116_ SKY130_FD_SC_HD__CLKINV_2
X_488_ NET176 VSSD VSSD VCCD VCCD _117_ SKY130_FD_SC_HD__CLKINV_2
X_489_ NET177 VSSD VSSD VCCD VCCD _118_ SKY130_FD_SC_HD__INV_2
X_490_ NET178 VSSD VSSD VCCD VCCD _119_ SKY130_FD_SC_HD__INV_2
X_491_ NET179 VSSD VSSD VCCD VCCD _120_ SKY130_FD_SC_HD__CLKINV_2
X_492_ NET180 VSSD VSSD VCCD VCCD _121_ SKY130_FD_SC_HD__CLKINV_2
X_493_ NET181 VSSD VSSD VCCD VCCD _122_ SKY130_FD_SC_HD__INV_2
X_494_ NET183 VSSD VSSD VCCD VCCD _124_ SKY130_FD_SC_HD__INV_2
X_495_ NET184 VSSD VSSD VCCD VCCD _125_ SKY130_FD_SC_HD__CLKINV_2
X_496_ NET185 VSSD VSSD VCCD VCCD _126_ SKY130_FD_SC_HD__INV_2
X_497_ NET186 VSSD VSSD VCCD VCCD _127_ SKY130_FD_SC_HD__CLKINV_2
X_498_ NET187 VSSD VSSD VCCD VCCD _128_ SKY130_FD_SC_HD__CLKINV_2
X_499_ NET188 VSSD VSSD VCCD VCCD _129_ SKY130_FD_SC_HD__CLKINV_2
X_500_ NET189 VSSD VSSD VCCD VCCD _130_ SKY130_FD_SC_HD__INV_2
X_501_ NET190 VSSD VSSD VCCD VCCD _131_ SKY130_FD_SC_HD__CLKINV_2
X_502_ NET191 VSSD VSSD VCCD VCCD _132_ SKY130_FD_SC_HD__CLKINV_2
X_503_ NET192 VSSD VSSD VCCD VCCD _133_ SKY130_FD_SC_HD__CLKINV_2
X_504_ NET194 VSSD VSSD VCCD VCCD _135_ SKY130_FD_SC_HD__CLKINV_2
X_505_ NET195 VSSD VSSD VCCD VCCD _136_ SKY130_FD_SC_HD__INV_2
X_506_ NET196 VSSD VSSD VCCD VCCD _137_ SKY130_FD_SC_HD__CLKINV_2
X_507_ NET197 VSSD VSSD VCCD VCCD _138_ SKY130_FD_SC_HD__CLKINV_2
X_508_ NET198 VSSD VSSD VCCD VCCD _139_ SKY130_FD_SC_HD__INV_2
X_509_ NET199 VSSD VSSD VCCD VCCD _140_ SKY130_FD_SC_HD__INV_2
X_510_ NET200 VSSD VSSD VCCD VCCD _141_ SKY130_FD_SC_HD__CLKINV_2
X_511_ NET201 VSSD VSSD VCCD VCCD _142_ SKY130_FD_SC_HD__CLKINV_2
X_512_ NET202 VSSD VSSD VCCD VCCD _143_ SKY130_FD_SC_HD__INV_2
X_513_ NET203 VSSD VSSD VCCD VCCD _144_ SKY130_FD_SC_HD__INV_2
X_514_ NET205 VSSD VSSD VCCD VCCD _146_ SKY130_FD_SC_HD__INV_2
X_515_ NET206 VSSD VSSD VCCD VCCD _147_ SKY130_FD_SC_HD__INV_2
X_516_ NET207 VSSD VSSD VCCD VCCD _148_ SKY130_FD_SC_HD__INV_2
X_517_ NET208 VSSD VSSD VCCD VCCD _149_ SKY130_FD_SC_HD__CLKINV_2
X_518_ NET209 VSSD VSSD VCCD VCCD _150_ SKY130_FD_SC_HD__INV_2
X_519_ NET210 VSSD VSSD VCCD VCCD _151_ SKY130_FD_SC_HD__CLKINV_2
X_520_ NET211 VSSD VSSD VCCD VCCD _152_ SKY130_FD_SC_HD__CLKINV_2
X_521_ NET212 VSSD VSSD VCCD VCCD _153_ SKY130_FD_SC_HD__INV_2
X_522_ NET213 VSSD VSSD VCCD VCCD _154_ SKY130_FD_SC_HD__INV_2
X_523_ NET214 VSSD VSSD VCCD VCCD _155_ SKY130_FD_SC_HD__CLKINV_2
X_524_ NET216 VSSD VSSD VCCD VCCD _157_ SKY130_FD_SC_HD__INV_2
X_525_ NET217 VSSD VSSD VCCD VCCD _158_ SKY130_FD_SC_HD__CLKINV_2
X_526_ NET218 VSSD VSSD VCCD VCCD _159_ SKY130_FD_SC_HD__CLKINV_2
X_527_ NET219 VSSD VSSD VCCD VCCD _160_ SKY130_FD_SC_HD__CLKINV_2
X_528_ NET220 VSSD VSSD VCCD VCCD _161_ SKY130_FD_SC_HD__CLKINV_2
X_529_ NET221 VSSD VSSD VCCD VCCD _162_ SKY130_FD_SC_HD__INV_2
X_530_ NET222 VSSD VSSD VCCD VCCD _163_ SKY130_FD_SC_HD__INV_2
X_531_ NET223 VSSD VSSD VCCD VCCD _164_ SKY130_FD_SC_HD__INV_2
X_532_ NET224 VSSD VSSD VCCD VCCD _165_ SKY130_FD_SC_HD__CLKINV_2
X_533_ NET225 VSSD VSSD VCCD VCCD _166_ SKY130_FD_SC_HD__INV_2
X_534_ NET227 VSSD VSSD VCCD VCCD _168_ SKY130_FD_SC_HD__CLKINV_2
X_535_ NET228 VSSD VSSD VCCD VCCD _169_ SKY130_FD_SC_HD__INV_2
X_536_ NET229 VSSD VSSD VCCD VCCD _170_ SKY130_FD_SC_HD__CLKINV_2
X_537_ NET230 VSSD VSSD VCCD VCCD _171_ SKY130_FD_SC_HD__INV_2
X_538_ NET231 VSSD VSSD VCCD VCCD _172_ SKY130_FD_SC_HD__CLKINV_2
X_539_ NET232 VSSD VSSD VCCD VCCD _173_ SKY130_FD_SC_HD__INV_2
X_540_ NET233 VSSD VSSD VCCD VCCD _174_ SKY130_FD_SC_HD__INV_2
X_541_ NET234 VSSD VSSD VCCD VCCD _175_ SKY130_FD_SC_HD__INV_2
X_542_ NET235 VSSD VSSD VCCD VCCD _176_ SKY130_FD_SC_HD__INV_2
X_543_ NET236 VSSD VSSD VCCD VCCD _177_ SKY130_FD_SC_HD__INV_2
X_544_ NET238 VSSD VSSD VCCD VCCD _179_ SKY130_FD_SC_HD__INV_2
X_545_ NET239 VSSD VSSD VCCD VCCD _180_ SKY130_FD_SC_HD__INV_2
X_546_ NET240 VSSD VSSD VCCD VCCD _181_ SKY130_FD_SC_HD__INV_2
X_547_ NET241 VSSD VSSD VCCD VCCD _182_ SKY130_FD_SC_HD__INV_2
X_548_ NET242 VSSD VSSD VCCD VCCD _183_ SKY130_FD_SC_HD__INV_2
X_549_ NET243 VSSD VSSD VCCD VCCD _184_ SKY130_FD_SC_HD__INV_2
X_550_ NET244 VSSD VSSD VCCD VCCD _185_ SKY130_FD_SC_HD__INV_2
X_551_ NET245 VSSD VSSD VCCD VCCD _186_ SKY130_FD_SC_HD__INV_2
X_552_ NET246 VSSD VSSD VCCD VCCD _187_ SKY130_FD_SC_HD__INV_2
X_553_ NET247 VSSD VSSD VCCD VCCD _188_ SKY130_FD_SC_HD__CLKINV_2
X_554_ NET249 VSSD VSSD VCCD VCCD _190_ SKY130_FD_SC_HD__INV_2
X_555_ NET250 VSSD VSSD VCCD VCCD _191_ SKY130_FD_SC_HD__CLKINV_2
X_556_ NET251 VSSD VSSD VCCD VCCD _192_ SKY130_FD_SC_HD__INV_2
X_557_ NET252 VSSD VSSD VCCD VCCD _193_ SKY130_FD_SC_HD__INV_2
X_558_ NET253 VSSD VSSD VCCD VCCD _194_ SKY130_FD_SC_HD__CLKINV_2
X_559_ NET254 VSSD VSSD VCCD VCCD _195_ SKY130_FD_SC_HD__INV_2
X_560_ NET255 VSSD VSSD VCCD VCCD _196_ SKY130_FD_SC_HD__INV_2
X_561_ NET256 VSSD VSSD VCCD VCCD _197_ SKY130_FD_SC_HD__INV_2
X_562_ NET257 VSSD VSSD VCCD VCCD _198_ SKY130_FD_SC_HD__CLKINV_2
X_563_ NET258 VSSD VSSD VCCD VCCD _199_ SKY130_FD_SC_HD__CLKINV_2
X_564_ NET133 VSSD VSSD VCCD VCCD _074_ SKY130_FD_SC_HD__CLKINV_2
X_565_ NET134 VSSD VSSD VCCD VCCD _075_ SKY130_FD_SC_HD__CLKINV_2
X_566_ NET135 VSSD VSSD VCCD VCCD _076_ SKY130_FD_SC_HD__INV_2
X_567_ NET136 VSSD VSSD VCCD VCCD _077_ SKY130_FD_SC_HD__INV_2
X_568_ NET137 VSSD VSSD VCCD VCCD _078_ SKY130_FD_SC_HD__CLKINV_2
X_569_ NET138 VSSD VSSD VCCD VCCD _079_ SKY130_FD_SC_HD__INV_2
X_570_ NET139 VSSD VSSD VCCD VCCD _080_ SKY130_FD_SC_HD__INV_2
X_571_ NET140 VSSD VSSD VCCD VCCD _081_ SKY130_FD_SC_HD__INV_2
X_572_ NET141 VSSD VSSD VCCD VCCD _082_ SKY130_FD_SC_HD__INV_2
X_573_ NET142 VSSD VSSD VCCD VCCD _083_ SKY130_FD_SC_HD__INV_2
X_574_ NET144 VSSD VSSD VCCD VCCD _085_ SKY130_FD_SC_HD__INV_2
X_575_ NET145 VSSD VSSD VCCD VCCD _086_ SKY130_FD_SC_HD__INV_2
X_576_ NET146 VSSD VSSD VCCD VCCD _087_ SKY130_FD_SC_HD__INV_2
X_577_ NET147 VSSD VSSD VCCD VCCD _088_ SKY130_FD_SC_HD__INV_2
X_578_ NET148 VSSD VSSD VCCD VCCD _089_ SKY130_FD_SC_HD__INV_2
X_579_ NET149 VSSD VSSD VCCD VCCD _090_ SKY130_FD_SC_HD__INV_2
X_580_ NET150 VSSD VSSD VCCD VCCD _091_ SKY130_FD_SC_HD__INV_2
X_581_ NET151 VSSD VSSD VCCD VCCD _092_ SKY130_FD_SC_HD__INV_2
X_582_ NET152 VSSD VSSD VCCD VCCD _093_ SKY130_FD_SC_HD__CLKINV_2
X_583_ NET153 VSSD VSSD VCCD VCCD _094_ SKY130_FD_SC_HD__INV_2
X_584_ NET155 VSSD VSSD VCCD VCCD _096_ SKY130_FD_SC_HD__CLKINV_2
X_585_ NET156 VSSD VSSD VCCD VCCD _097_ SKY130_FD_SC_HD__INV_2
X_586_ NET157 VSSD VSSD VCCD VCCD _098_ SKY130_FD_SC_HD__CLKINV_2
X_587_ NET158 VSSD VSSD VCCD VCCD _099_ SKY130_FD_SC_HD__INV_2
X_588_ NET159 VSSD VSSD VCCD VCCD _100_ SKY130_FD_SC_HD__INV_2
X_589_ NET160 VSSD VSSD VCCD VCCD _101_ SKY130_FD_SC_HD__CLKINV_2
X_590_ NET161 VSSD VSSD VCCD VCCD _102_ SKY130_FD_SC_HD__INV_2
X_591_ NET162 VSSD VSSD VCCD VCCD _103_ SKY130_FD_SC_HD__INV_2
X_592_ NET388 VSSD VSSD VCCD VCCD _201_ SKY130_FD_SC_HD__INV_2
X_593_ NET427 VSSD VSSD VCCD VCCD _240_ SKY130_FD_SC_HD__INV_2
X_594_ NET438 VSSD VSSD VCCD VCCD _251_ SKY130_FD_SC_HD__CLKINV_2
X_595_ NET449 VSSD VSSD VCCD VCCD _262_ SKY130_FD_SC_HD__INV_2
X_596_ NET460 VSSD VSSD VCCD VCCD _273_ SKY130_FD_SC_HD__INV_2
X_597_ NET471 VSSD VSSD VCCD VCCD _284_ SKY130_FD_SC_HD__CLKINV_2
X_598_ NET482 VSSD VSSD VCCD VCCD _295_ SKY130_FD_SC_HD__INV_2
X_599_ NET493 VSSD VSSD VCCD VCCD _306_ SKY130_FD_SC_HD__INV_2
X_600_ NET504 VSSD VSSD VCCD VCCD _317_ SKY130_FD_SC_HD__CLKINV_2
X_601_ NET515 VSSD VSSD VCCD VCCD _328_ SKY130_FD_SC_HD__INV_2
X_602_ NET399 VSSD VSSD VCCD VCCD _212_ SKY130_FD_SC_HD__INV_2
X_603_ NET410 VSSD VSSD VCCD VCCD _223_ SKY130_FD_SC_HD__INV_2
X_604_ NET419 VSSD VSSD VCCD VCCD _232_ SKY130_FD_SC_HD__CLKINV_2
X_605_ NET420 VSSD VSSD VCCD VCCD _233_ SKY130_FD_SC_HD__INV_2
X_606_ NET421 VSSD VSSD VCCD VCCD _234_ SKY130_FD_SC_HD__CLKINV_2
X_607_ NET422 VSSD VSSD VCCD VCCD _235_ SKY130_FD_SC_HD__CLKINV_2
X_608_ NET423 VSSD VSSD VCCD VCCD _236_ SKY130_FD_SC_HD__INV_2
X_609_ NET424 VSSD VSSD VCCD VCCD _237_ SKY130_FD_SC_HD__CLKINV_2
X_610_ NET425 VSSD VSSD VCCD VCCD _238_ SKY130_FD_SC_HD__INV_2
X_611_ NET426 VSSD VSSD VCCD VCCD _239_ SKY130_FD_SC_HD__CLKINV_2
X_612_ NET428 VSSD VSSD VCCD VCCD _241_ SKY130_FD_SC_HD__INV_2
X_613_ NET429 VSSD VSSD VCCD VCCD _242_ SKY130_FD_SC_HD__INV_2
X_614_ NET430 VSSD VSSD VCCD VCCD _243_ SKY130_FD_SC_HD__INV_2
X_615_ NET431 VSSD VSSD VCCD VCCD _244_ SKY130_FD_SC_HD__INV_2
X_616_ NET432 VSSD VSSD VCCD VCCD _245_ SKY130_FD_SC_HD__CLKINV_2
X_617_ NET433 VSSD VSSD VCCD VCCD _246_ SKY130_FD_SC_HD__CLKINV_2
X_618_ NET434 VSSD VSSD VCCD VCCD _247_ SKY130_FD_SC_HD__CLKINV_2
X_619_ NET435 VSSD VSSD VCCD VCCD _248_ SKY130_FD_SC_HD__CLKINV_2
X_620_ NET436 VSSD VSSD VCCD VCCD _249_ SKY130_FD_SC_HD__CLKINV_2
X_621_ NET437 VSSD VSSD VCCD VCCD _250_ SKY130_FD_SC_HD__CLKINV_2
X_622_ NET439 VSSD VSSD VCCD VCCD _252_ SKY130_FD_SC_HD__INV_2
X_623_ NET440 VSSD VSSD VCCD VCCD _253_ SKY130_FD_SC_HD__CLKINV_2
X_624_ NET441 VSSD VSSD VCCD VCCD _254_ SKY130_FD_SC_HD__CLKINV_2
X_625_ NET442 VSSD VSSD VCCD VCCD _255_ SKY130_FD_SC_HD__CLKINV_2
X_626_ NET443 VSSD VSSD VCCD VCCD _256_ SKY130_FD_SC_HD__INV_2
X_627_ NET444 VSSD VSSD VCCD VCCD _257_ SKY130_FD_SC_HD__INV_2
X_628_ NET445 VSSD VSSD VCCD VCCD _258_ SKY130_FD_SC_HD__INV_2
X_629_ NET446 VSSD VSSD VCCD VCCD _259_ SKY130_FD_SC_HD__INV_2
X_630_ NET447 VSSD VSSD VCCD VCCD _260_ SKY130_FD_SC_HD__INV_2
X_631_ NET448 VSSD VSSD VCCD VCCD _261_ SKY130_FD_SC_HD__INV_2
X_632_ NET450 VSSD VSSD VCCD VCCD _263_ SKY130_FD_SC_HD__INV_2
X_633_ NET451 VSSD VSSD VCCD VCCD _264_ SKY130_FD_SC_HD__CLKINV_2
X_634_ NET452 VSSD VSSD VCCD VCCD _265_ SKY130_FD_SC_HD__INV_2
X_635_ NET453 VSSD VSSD VCCD VCCD _266_ SKY130_FD_SC_HD__INV_2
X_636_ NET454 VSSD VSSD VCCD VCCD _267_ SKY130_FD_SC_HD__INV_2
X_637_ NET455 VSSD VSSD VCCD VCCD _268_ SKY130_FD_SC_HD__CLKINV_2
X_638_ NET456 VSSD VSSD VCCD VCCD _269_ SKY130_FD_SC_HD__INV_2
X_639_ NET457 VSSD VSSD VCCD VCCD _270_ SKY130_FD_SC_HD__INV_2
X_640_ NET458 VSSD VSSD VCCD VCCD _271_ SKY130_FD_SC_HD__INV_2
X_641_ NET459 VSSD VSSD VCCD VCCD _272_ SKY130_FD_SC_HD__INV_2
X_642_ NET461 VSSD VSSD VCCD VCCD _274_ SKY130_FD_SC_HD__CLKINV_2
X_643_ NET462 VSSD VSSD VCCD VCCD _275_ SKY130_FD_SC_HD__INV_2
X_644_ NET463 VSSD VSSD VCCD VCCD _276_ SKY130_FD_SC_HD__CLKINV_2
X_645_ NET464 VSSD VSSD VCCD VCCD _277_ SKY130_FD_SC_HD__CLKINV_2
X_646_ NET465 VSSD VSSD VCCD VCCD _278_ SKY130_FD_SC_HD__INV_2
X_647_ NET466 VSSD VSSD VCCD VCCD _279_ SKY130_FD_SC_HD__CLKINV_2
X_648_ NET467 VSSD VSSD VCCD VCCD _280_ SKY130_FD_SC_HD__CLKINV_2
X_649_ NET468 VSSD VSSD VCCD VCCD _281_ SKY130_FD_SC_HD__CLKINV_2
X_650_ NET469 VSSD VSSD VCCD VCCD _282_ SKY130_FD_SC_HD__CLKINV_2
X_651_ NET470 VSSD VSSD VCCD VCCD _283_ SKY130_FD_SC_HD__CLKINV_2
X_652_ NET472 VSSD VSSD VCCD VCCD _285_ SKY130_FD_SC_HD__INV_2
X_653_ NET473 VSSD VSSD VCCD VCCD _286_ SKY130_FD_SC_HD__INV_2
X_654_ NET474 VSSD VSSD VCCD VCCD _287_ SKY130_FD_SC_HD__INV_2
X_655_ NET475 VSSD VSSD VCCD VCCD _288_ SKY130_FD_SC_HD__CLKINV_2
X_656_ NET476 VSSD VSSD VCCD VCCD _289_ SKY130_FD_SC_HD__INV_2
X_657_ NET477 VSSD VSSD VCCD VCCD _290_ SKY130_FD_SC_HD__INV_2
XINPUT1 CARAVEL_CLK VSSD VSSD VCCD VCCD NET1 SKY130_FD_SC_HD__CLKBUF_1
XINPUT10 LA_DATA_OUT_CORE[105] VSSD VSSD VCCD VCCD NET10 SKY130_FD_SC_HD__BUF_4
XINPUT100 LA_DATA_OUT_CORE[71] VSSD VSSD VCCD VCCD NET100 SKY130_FD_SC_HD__BUF_4
XINPUT101 LA_DATA_OUT_CORE[72] VSSD VSSD VCCD VCCD NET101 SKY130_FD_SC_HD__BUF_4
XINPUT102 LA_DATA_OUT_CORE[73] VSSD VSSD VCCD VCCD NET102 SKY130_FD_SC_HD__BUF_4
XINPUT103 LA_DATA_OUT_CORE[74] VSSD VSSD VCCD VCCD NET103 SKY130_FD_SC_HD__BUF_4
XINPUT104 LA_DATA_OUT_CORE[75] VSSD VSSD VCCD VCCD NET104 SKY130_FD_SC_HD__BUF_4
XINPUT105 LA_DATA_OUT_CORE[76] VSSD VSSD VCCD VCCD NET105 SKY130_FD_SC_HD__BUF_4
XINPUT106 LA_DATA_OUT_CORE[77] VSSD VSSD VCCD VCCD NET106 SKY130_FD_SC_HD__BUF_4
XINPUT107 LA_DATA_OUT_CORE[78] VSSD VSSD VCCD VCCD NET107 SKY130_FD_SC_HD__BUF_4
XINPUT108 LA_DATA_OUT_CORE[79] VSSD VSSD VCCD VCCD NET108 SKY130_FD_SC_HD__BUF_4
XINPUT109 LA_DATA_OUT_CORE[7] VSSD VSSD VCCD VCCD NET109 SKY130_FD_SC_HD__CLKBUF_4
XINPUT11 LA_DATA_OUT_CORE[106] VSSD VSSD VCCD VCCD NET11 SKY130_FD_SC_HD__BUF_4
XINPUT110 LA_DATA_OUT_CORE[80] VSSD VSSD VCCD VCCD NET110 SKY130_FD_SC_HD__BUF_4
XINPUT111 LA_DATA_OUT_CORE[81] VSSD VSSD VCCD VCCD NET111 SKY130_FD_SC_HD__BUF_4
XINPUT112 LA_DATA_OUT_CORE[82] VSSD VSSD VCCD VCCD NET112 SKY130_FD_SC_HD__BUF_4
XINPUT113 LA_DATA_OUT_CORE[83] VSSD VSSD VCCD VCCD NET113 SKY130_FD_SC_HD__BUF_4
XINPUT114 LA_DATA_OUT_CORE[84] VSSD VSSD VCCD VCCD NET114 SKY130_FD_SC_HD__BUF_4
XINPUT115 LA_DATA_OUT_CORE[85] VSSD VSSD VCCD VCCD NET115 SKY130_FD_SC_HD__BUF_4
XINPUT116 LA_DATA_OUT_CORE[86] VSSD VSSD VCCD VCCD NET116 SKY130_FD_SC_HD__BUF_4
XINPUT117 LA_DATA_OUT_CORE[87] VSSD VSSD VCCD VCCD NET117 SKY130_FD_SC_HD__BUF_4
XINPUT118 LA_DATA_OUT_CORE[88] VSSD VSSD VCCD VCCD NET118 SKY130_FD_SC_HD__BUF_4
XINPUT119 LA_DATA_OUT_CORE[89] VSSD VSSD VCCD VCCD NET119 SKY130_FD_SC_HD__BUF_4
XINPUT12 LA_DATA_OUT_CORE[107] VSSD VSSD VCCD VCCD NET12 SKY130_FD_SC_HD__BUF_4
XINPUT120 LA_DATA_OUT_CORE[8] VSSD VSSD VCCD VCCD NET120 SKY130_FD_SC_HD__CLKBUF_4
XINPUT121 LA_DATA_OUT_CORE[90] VSSD VSSD VCCD VCCD NET121 SKY130_FD_SC_HD__BUF_4
XINPUT122 LA_DATA_OUT_CORE[91] VSSD VSSD VCCD VCCD NET122 SKY130_FD_SC_HD__CLKBUF_4
XINPUT123 LA_DATA_OUT_CORE[92] VSSD VSSD VCCD VCCD NET123 SKY130_FD_SC_HD__BUF_4
XINPUT124 LA_DATA_OUT_CORE[93] VSSD VSSD VCCD VCCD NET124 SKY130_FD_SC_HD__BUF_4
XINPUT125 LA_DATA_OUT_CORE[94] VSSD VSSD VCCD VCCD NET125 SKY130_FD_SC_HD__BUF_4
XINPUT126 LA_DATA_OUT_CORE[95] VSSD VSSD VCCD VCCD NET126 SKY130_FD_SC_HD__BUF_4
XINPUT127 LA_DATA_OUT_CORE[96] VSSD VSSD VCCD VCCD NET127 SKY130_FD_SC_HD__BUF_4
XINPUT128 LA_DATA_OUT_CORE[97] VSSD VSSD VCCD VCCD NET128 SKY130_FD_SC_HD__BUF_4
XINPUT129 LA_DATA_OUT_CORE[98] VSSD VSSD VCCD VCCD NET129 SKY130_FD_SC_HD__BUF_4
XINPUT13 LA_DATA_OUT_CORE[108] VSSD VSSD VCCD VCCD NET13 SKY130_FD_SC_HD__CLKBUF_4
XINPUT130 LA_DATA_OUT_CORE[99] VSSD VSSD VCCD VCCD NET130 SKY130_FD_SC_HD__CLKBUF_4
XINPUT131 LA_DATA_OUT_CORE[9] VSSD VSSD VCCD VCCD NET131 SKY130_FD_SC_HD__BUF_2
XINPUT132 LA_DATA_OUT_MPRJ[0] VSSD VSSD VCCD VCCD NET132 SKY130_FD_SC_HD__CLKBUF_2
XINPUT133 LA_DATA_OUT_MPRJ[100] VSSD VSSD VCCD VCCD NET133 SKY130_FD_SC_HD__BUF_2
XINPUT134 LA_DATA_OUT_MPRJ[101] VSSD VSSD VCCD VCCD NET134 SKY130_FD_SC_HD__BUF_2
XINPUT135 LA_DATA_OUT_MPRJ[102] VSSD VSSD VCCD VCCD NET135 SKY130_FD_SC_HD__CLKBUF_4
XINPUT136 LA_DATA_OUT_MPRJ[103] VSSD VSSD VCCD VCCD NET136 SKY130_FD_SC_HD__CLKBUF_4
XINPUT137 LA_DATA_OUT_MPRJ[104] VSSD VSSD VCCD VCCD NET137 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT138 LA_DATA_OUT_MPRJ[105] VSSD VSSD VCCD VCCD NET138 SKY130_FD_SC_HD__CLKBUF_2
XINPUT139 LA_DATA_OUT_MPRJ[106] VSSD VSSD VCCD VCCD NET139 SKY130_FD_SC_HD__CLKBUF_2
XINPUT14 LA_DATA_OUT_CORE[109] VSSD VSSD VCCD VCCD NET14 SKY130_FD_SC_HD__CLKBUF_4
XINPUT140 LA_DATA_OUT_MPRJ[107] VSSD VSSD VCCD VCCD NET140 SKY130_FD_SC_HD__CLKBUF_4
XINPUT141 LA_DATA_OUT_MPRJ[108] VSSD VSSD VCCD VCCD NET141 SKY130_FD_SC_HD__CLKBUF_2
XINPUT142 LA_DATA_OUT_MPRJ[109] VSSD VSSD VCCD VCCD NET142 SKY130_FD_SC_HD__CLKBUF_4
XINPUT143 LA_DATA_OUT_MPRJ[10] VSSD VSSD VCCD VCCD NET143 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT144 LA_DATA_OUT_MPRJ[110] VSSD VSSD VCCD VCCD NET144 SKY130_FD_SC_HD__CLKBUF_4
XINPUT145 LA_DATA_OUT_MPRJ[111] VSSD VSSD VCCD VCCD NET145 SKY130_FD_SC_HD__CLKBUF_4
XINPUT146 LA_DATA_OUT_MPRJ[112] VSSD VSSD VCCD VCCD NET146 SKY130_FD_SC_HD__CLKBUF_4
XINPUT147 LA_DATA_OUT_MPRJ[113] VSSD VSSD VCCD VCCD NET147 SKY130_FD_SC_HD__CLKBUF_4
XINPUT148 LA_DATA_OUT_MPRJ[114] VSSD VSSD VCCD VCCD NET148 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT149 LA_DATA_OUT_MPRJ[115] VSSD VSSD VCCD VCCD NET149 SKY130_FD_SC_HD__BUF_2
XINPUT15 LA_DATA_OUT_CORE[10] VSSD VSSD VCCD VCCD NET15 SKY130_FD_SC_HD__BUF_2
XINPUT150 LA_DATA_OUT_MPRJ[116] VSSD VSSD VCCD VCCD NET150 SKY130_FD_SC_HD__CLKBUF_2
XINPUT151 LA_DATA_OUT_MPRJ[117] VSSD VSSD VCCD VCCD NET151 SKY130_FD_SC_HD__CLKBUF_4
XINPUT152 LA_DATA_OUT_MPRJ[118] VSSD VSSD VCCD VCCD NET152 SKY130_FD_SC_HD__CLKBUF_2
XINPUT153 LA_DATA_OUT_MPRJ[119] VSSD VSSD VCCD VCCD NET153 SKY130_FD_SC_HD__CLKBUF_4
XINPUT154 LA_DATA_OUT_MPRJ[11] VSSD VSSD VCCD VCCD NET154 SKY130_FD_SC_HD__CLKBUF_2
XINPUT155 LA_DATA_OUT_MPRJ[120] VSSD VSSD VCCD VCCD NET155 SKY130_FD_SC_HD__CLKBUF_2
XINPUT156 LA_DATA_OUT_MPRJ[121] VSSD VSSD VCCD VCCD NET156 SKY130_FD_SC_HD__CLKBUF_2
XINPUT157 LA_DATA_OUT_MPRJ[122] VSSD VSSD VCCD VCCD NET157 SKY130_FD_SC_HD__CLKBUF_2
XINPUT158 LA_DATA_OUT_MPRJ[123] VSSD VSSD VCCD VCCD NET158 SKY130_FD_SC_HD__CLKBUF_4
XINPUT159 LA_DATA_OUT_MPRJ[124] VSSD VSSD VCCD VCCD NET159 SKY130_FD_SC_HD__CLKBUF_4
XINPUT16 LA_DATA_OUT_CORE[110] VSSD VSSD VCCD VCCD NET16 SKY130_FD_SC_HD__BUF_4
XINPUT160 LA_DATA_OUT_MPRJ[125] VSSD VSSD VCCD VCCD NET160 SKY130_FD_SC_HD__CLKBUF_2
XINPUT161 LA_DATA_OUT_MPRJ[126] VSSD VSSD VCCD VCCD NET161 SKY130_FD_SC_HD__CLKBUF_4
XINPUT162 LA_DATA_OUT_MPRJ[127] VSSD VSSD VCCD VCCD NET162 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT163 LA_DATA_OUT_MPRJ[12] VSSD VSSD VCCD VCCD NET163 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT164 LA_DATA_OUT_MPRJ[13] VSSD VSSD VCCD VCCD NET164 SKY130_FD_SC_HD__CLKBUF_2
XINPUT165 LA_DATA_OUT_MPRJ[14] VSSD VSSD VCCD VCCD NET165 SKY130_FD_SC_HD__CLKBUF_2
XINPUT166 LA_DATA_OUT_MPRJ[15] VSSD VSSD VCCD VCCD NET166 SKY130_FD_SC_HD__CLKBUF_2
XINPUT167 LA_DATA_OUT_MPRJ[16] VSSD VSSD VCCD VCCD NET167 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT168 LA_DATA_OUT_MPRJ[17] VSSD VSSD VCCD VCCD NET168 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT169 LA_DATA_OUT_MPRJ[18] VSSD VSSD VCCD VCCD NET169 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT17 LA_DATA_OUT_CORE[111] VSSD VSSD VCCD VCCD NET17 SKY130_FD_SC_HD__BUF_4
XINPUT170 LA_DATA_OUT_MPRJ[19] VSSD VSSD VCCD VCCD NET170 SKY130_FD_SC_HD__CLKBUF_2
XINPUT171 LA_DATA_OUT_MPRJ[1] VSSD VSSD VCCD VCCD NET171 SKY130_FD_SC_HD__CLKBUF_2
XINPUT172 LA_DATA_OUT_MPRJ[20] VSSD VSSD VCCD VCCD NET172 SKY130_FD_SC_HD__CLKBUF_2
XINPUT173 LA_DATA_OUT_MPRJ[21] VSSD VSSD VCCD VCCD NET173 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT174 LA_DATA_OUT_MPRJ[22] VSSD VSSD VCCD VCCD NET174 SKY130_FD_SC_HD__CLKBUF_2
XINPUT175 LA_DATA_OUT_MPRJ[23] VSSD VSSD VCCD VCCD NET175 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT176 LA_DATA_OUT_MPRJ[24] VSSD VSSD VCCD VCCD NET176 SKY130_FD_SC_HD__CLKBUF_2
XINPUT177 LA_DATA_OUT_MPRJ[25] VSSD VSSD VCCD VCCD NET177 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT178 LA_DATA_OUT_MPRJ[26] VSSD VSSD VCCD VCCD NET178 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT179 LA_DATA_OUT_MPRJ[27] VSSD VSSD VCCD VCCD NET179 SKY130_FD_SC_HD__CLKBUF_2
XINPUT18 LA_DATA_OUT_CORE[112] VSSD VSSD VCCD VCCD NET18 SKY130_FD_SC_HD__CLKBUF_4
XINPUT180 LA_DATA_OUT_MPRJ[28] VSSD VSSD VCCD VCCD NET180 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT181 LA_DATA_OUT_MPRJ[29] VSSD VSSD VCCD VCCD NET181 SKY130_FD_SC_HD__CLKBUF_2
XINPUT182 LA_DATA_OUT_MPRJ[2] VSSD VSSD VCCD VCCD NET182 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT183 LA_DATA_OUT_MPRJ[30] VSSD VSSD VCCD VCCD NET183 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT184 LA_DATA_OUT_MPRJ[31] VSSD VSSD VCCD VCCD NET184 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT185 LA_DATA_OUT_MPRJ[32] VSSD VSSD VCCD VCCD NET185 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT186 LA_DATA_OUT_MPRJ[33] VSSD VSSD VCCD VCCD NET186 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT187 LA_DATA_OUT_MPRJ[34] VSSD VSSD VCCD VCCD NET187 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT188 LA_DATA_OUT_MPRJ[35] VSSD VSSD VCCD VCCD NET188 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT189 LA_DATA_OUT_MPRJ[36] VSSD VSSD VCCD VCCD NET189 SKY130_FD_SC_HD__CLKBUF_1
XINPUT19 LA_DATA_OUT_CORE[113] VSSD VSSD VCCD VCCD NET19 SKY130_FD_SC_HD__CLKBUF_4
XINPUT190 LA_DATA_OUT_MPRJ[37] VSSD VSSD VCCD VCCD NET190 SKY130_FD_SC_HD__CLKBUF_1
XINPUT191 LA_DATA_OUT_MPRJ[38] VSSD VSSD VCCD VCCD NET191 SKY130_FD_SC_HD__CLKBUF_1
XINPUT192 LA_DATA_OUT_MPRJ[39] VSSD VSSD VCCD VCCD NET192 SKY130_FD_SC_HD__CLKBUF_1
XINPUT193 LA_DATA_OUT_MPRJ[3] VSSD VSSD VCCD VCCD NET193 SKY130_FD_SC_HD__CLKBUF_2
XINPUT194 LA_DATA_OUT_MPRJ[40] VSSD VSSD VCCD VCCD NET194 SKY130_FD_SC_HD__CLKBUF_2
XINPUT195 LA_DATA_OUT_MPRJ[41] VSSD VSSD VCCD VCCD NET195 SKY130_FD_SC_HD__CLKBUF_2
XINPUT196 LA_DATA_OUT_MPRJ[42] VSSD VSSD VCCD VCCD NET196 SKY130_FD_SC_HD__CLKBUF_2
XINPUT197 LA_DATA_OUT_MPRJ[43] VSSD VSSD VCCD VCCD NET197 SKY130_FD_SC_HD__CLKBUF_2
XINPUT198 LA_DATA_OUT_MPRJ[44] VSSD VSSD VCCD VCCD NET198 SKY130_FD_SC_HD__CLKBUF_2
XINPUT199 LA_DATA_OUT_MPRJ[45] VSSD VSSD VCCD VCCD NET199 SKY130_FD_SC_HD__CLKBUF_2
XINPUT2 CARAVEL_CLK2 VSSD VSSD VCCD VCCD NET2 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT20 LA_DATA_OUT_CORE[114] VSSD VSSD VCCD VCCD NET20 SKY130_FD_SC_HD__CLKBUF_4
XINPUT200 LA_DATA_OUT_MPRJ[46] VSSD VSSD VCCD VCCD NET200 SKY130_FD_SC_HD__CLKBUF_2
XINPUT201 LA_DATA_OUT_MPRJ[47] VSSD VSSD VCCD VCCD NET201 SKY130_FD_SC_HD__CLKBUF_2
XINPUT202 LA_DATA_OUT_MPRJ[48] VSSD VSSD VCCD VCCD NET202 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT203 LA_DATA_OUT_MPRJ[49] VSSD VSSD VCCD VCCD NET203 SKY130_FD_SC_HD__CLKBUF_2
XINPUT204 LA_DATA_OUT_MPRJ[4] VSSD VSSD VCCD VCCD NET204 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT205 LA_DATA_OUT_MPRJ[50] VSSD VSSD VCCD VCCD NET205 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT206 LA_DATA_OUT_MPRJ[51] VSSD VSSD VCCD VCCD NET206 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT207 LA_DATA_OUT_MPRJ[52] VSSD VSSD VCCD VCCD NET207 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT208 LA_DATA_OUT_MPRJ[53] VSSD VSSD VCCD VCCD NET208 SKY130_FD_SC_HD__CLKBUF_2
XINPUT209 LA_DATA_OUT_MPRJ[54] VSSD VSSD VCCD VCCD NET209 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT21 LA_DATA_OUT_CORE[115] VSSD VSSD VCCD VCCD NET21 SKY130_FD_SC_HD__CLKBUF_4
XINPUT210 LA_DATA_OUT_MPRJ[55] VSSD VSSD VCCD VCCD NET210 SKY130_FD_SC_HD__CLKBUF_2
XINPUT211 LA_DATA_OUT_MPRJ[56] VSSD VSSD VCCD VCCD NET211 SKY130_FD_SC_HD__CLKBUF_2
XINPUT212 LA_DATA_OUT_MPRJ[57] VSSD VSSD VCCD VCCD NET212 SKY130_FD_SC_HD__CLKBUF_2
XINPUT213 LA_DATA_OUT_MPRJ[58] VSSD VSSD VCCD VCCD NET213 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT214 LA_DATA_OUT_MPRJ[59] VSSD VSSD VCCD VCCD NET214 SKY130_FD_SC_HD__CLKBUF_2
XINPUT215 LA_DATA_OUT_MPRJ[5] VSSD VSSD VCCD VCCD NET215 SKY130_FD_SC_HD__CLKBUF_2
XINPUT216 LA_DATA_OUT_MPRJ[60] VSSD VSSD VCCD VCCD NET216 SKY130_FD_SC_HD__CLKBUF_2
XINPUT217 LA_DATA_OUT_MPRJ[61] VSSD VSSD VCCD VCCD NET217 SKY130_FD_SC_HD__CLKBUF_2
XINPUT218 LA_DATA_OUT_MPRJ[62] VSSD VSSD VCCD VCCD NET218 SKY130_FD_SC_HD__CLKBUF_2
XINPUT219 LA_DATA_OUT_MPRJ[63] VSSD VSSD VCCD VCCD NET219 SKY130_FD_SC_HD__CLKBUF_2
XINPUT22 LA_DATA_OUT_CORE[116] VSSD VSSD VCCD VCCD NET22 SKY130_FD_SC_HD__CLKBUF_4
XINPUT220 LA_DATA_OUT_MPRJ[64] VSSD VSSD VCCD VCCD NET220 SKY130_FD_SC_HD__BUF_2
XINPUT221 LA_DATA_OUT_MPRJ[65] VSSD VSSD VCCD VCCD NET221 SKY130_FD_SC_HD__CLKBUF_2
XINPUT222 LA_DATA_OUT_MPRJ[66] VSSD VSSD VCCD VCCD NET222 SKY130_FD_SC_HD__CLKBUF_2
XINPUT223 LA_DATA_OUT_MPRJ[67] VSSD VSSD VCCD VCCD NET223 SKY130_FD_SC_HD__CLKBUF_2
XINPUT224 LA_DATA_OUT_MPRJ[68] VSSD VSSD VCCD VCCD NET224 SKY130_FD_SC_HD__CLKBUF_2
XINPUT225 LA_DATA_OUT_MPRJ[69] VSSD VSSD VCCD VCCD NET225 SKY130_FD_SC_HD__CLKBUF_2
XINPUT226 LA_DATA_OUT_MPRJ[6] VSSD VSSD VCCD VCCD NET226 SKY130_FD_SC_HD__CLKBUF_2
XINPUT227 LA_DATA_OUT_MPRJ[70] VSSD VSSD VCCD VCCD NET227 SKY130_FD_SC_HD__BUF_2
XINPUT228 LA_DATA_OUT_MPRJ[71] VSSD VSSD VCCD VCCD NET228 SKY130_FD_SC_HD__BUF_2
XINPUT229 LA_DATA_OUT_MPRJ[72] VSSD VSSD VCCD VCCD NET229 SKY130_FD_SC_HD__CLKBUF_2
XINPUT23 LA_DATA_OUT_CORE[117] VSSD VSSD VCCD VCCD NET23 SKY130_FD_SC_HD__BUF_4
XINPUT230 LA_DATA_OUT_MPRJ[73] VSSD VSSD VCCD VCCD NET230 SKY130_FD_SC_HD__BUF_2
XINPUT231 LA_DATA_OUT_MPRJ[74] VSSD VSSD VCCD VCCD NET231 SKY130_FD_SC_HD__CLKBUF_2
XINPUT232 LA_DATA_OUT_MPRJ[75] VSSD VSSD VCCD VCCD NET232 SKY130_FD_SC_HD__BUF_2
XINPUT233 LA_DATA_OUT_MPRJ[76] VSSD VSSD VCCD VCCD NET233 SKY130_FD_SC_HD__CLKBUF_4
XINPUT234 LA_DATA_OUT_MPRJ[77] VSSD VSSD VCCD VCCD NET234 SKY130_FD_SC_HD__BUF_2
XINPUT235 LA_DATA_OUT_MPRJ[78] VSSD VSSD VCCD VCCD NET235 SKY130_FD_SC_HD__CLKBUF_4
XINPUT236 LA_DATA_OUT_MPRJ[79] VSSD VSSD VCCD VCCD NET236 SKY130_FD_SC_HD__CLKBUF_4
XINPUT237 LA_DATA_OUT_MPRJ[7] VSSD VSSD VCCD VCCD NET237 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT238 LA_DATA_OUT_MPRJ[80] VSSD VSSD VCCD VCCD NET238 SKY130_FD_SC_HD__BUF_4
XINPUT239 LA_DATA_OUT_MPRJ[81] VSSD VSSD VCCD VCCD NET239 SKY130_FD_SC_HD__CLKBUF_4
XINPUT24 LA_DATA_OUT_CORE[118] VSSD VSSD VCCD VCCD NET24 SKY130_FD_SC_HD__CLKBUF_4
XINPUT240 LA_DATA_OUT_MPRJ[82] VSSD VSSD VCCD VCCD NET240 SKY130_FD_SC_HD__BUF_4
XINPUT241 LA_DATA_OUT_MPRJ[83] VSSD VSSD VCCD VCCD NET241 SKY130_FD_SC_HD__BUF_4
XINPUT242 LA_DATA_OUT_MPRJ[84] VSSD VSSD VCCD VCCD NET242 SKY130_FD_SC_HD__BUF_4
XINPUT243 LA_DATA_OUT_MPRJ[85] VSSD VSSD VCCD VCCD NET243 SKY130_FD_SC_HD__BUF_4
XINPUT244 LA_DATA_OUT_MPRJ[86] VSSD VSSD VCCD VCCD NET244 SKY130_FD_SC_HD__CLKBUF_4
XINPUT245 LA_DATA_OUT_MPRJ[87] VSSD VSSD VCCD VCCD NET245 SKY130_FD_SC_HD__BUF_2
XINPUT246 LA_DATA_OUT_MPRJ[88] VSSD VSSD VCCD VCCD NET246 SKY130_FD_SC_HD__CLKBUF_4
XINPUT247 LA_DATA_OUT_MPRJ[89] VSSD VSSD VCCD VCCD NET247 SKY130_FD_SC_HD__CLKBUF_1
XINPUT248 LA_DATA_OUT_MPRJ[8] VSSD VSSD VCCD VCCD NET248 SKY130_FD_SC_HD__CLKBUF_2
XINPUT249 LA_DATA_OUT_MPRJ[90] VSSD VSSD VCCD VCCD NET249 SKY130_FD_SC_HD__CLKBUF_2
XINPUT25 LA_DATA_OUT_CORE[119] VSSD VSSD VCCD VCCD NET25 SKY130_FD_SC_HD__BUF_2
XINPUT250 LA_DATA_OUT_MPRJ[91] VSSD VSSD VCCD VCCD NET250 SKY130_FD_SC_HD__CLKBUF_1
XINPUT251 LA_DATA_OUT_MPRJ[92] VSSD VSSD VCCD VCCD NET251 SKY130_FD_SC_HD__CLKBUF_2
XINPUT252 LA_DATA_OUT_MPRJ[93] VSSD VSSD VCCD VCCD NET252 SKY130_FD_SC_HD__BUF_2
XINPUT253 LA_DATA_OUT_MPRJ[94] VSSD VSSD VCCD VCCD NET253 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT254 LA_DATA_OUT_MPRJ[95] VSSD VSSD VCCD VCCD NET254 SKY130_FD_SC_HD__CLKBUF_2
XINPUT255 LA_DATA_OUT_MPRJ[96] VSSD VSSD VCCD VCCD NET255 SKY130_FD_SC_HD__BUF_2
XINPUT256 LA_DATA_OUT_MPRJ[97] VSSD VSSD VCCD VCCD NET256 SKY130_FD_SC_HD__BUF_2
XINPUT257 LA_DATA_OUT_MPRJ[98] VSSD VSSD VCCD VCCD NET257 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT258 LA_DATA_OUT_MPRJ[99] VSSD VSSD VCCD VCCD NET258 SKY130_FD_SC_HD__CLKBUF_1
XINPUT259 LA_DATA_OUT_MPRJ[9] VSSD VSSD VCCD VCCD NET259 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT26 LA_DATA_OUT_CORE[11] VSSD VSSD VCCD VCCD NET26 SKY130_FD_SC_HD__CLKBUF_4
XINPUT260 LA_IENA_MPRJ[0] VSSD VSSD VCCD VCCD NET260 SKY130_FD_SC_HD__CLKBUF_1
XINPUT261 LA_IENA_MPRJ[100] VSSD VSSD VCCD VCCD NET261 SKY130_FD_SC_HD__CLKBUF_1
XINPUT262 LA_IENA_MPRJ[101] VSSD VSSD VCCD VCCD NET262 SKY130_FD_SC_HD__CLKBUF_1
XINPUT263 LA_IENA_MPRJ[102] VSSD VSSD VCCD VCCD NET263 SKY130_FD_SC_HD__CLKBUF_1
XINPUT264 LA_IENA_MPRJ[103] VSSD VSSD VCCD VCCD NET264 SKY130_FD_SC_HD__CLKBUF_1
XINPUT265 LA_IENA_MPRJ[104] VSSD VSSD VCCD VCCD NET265 SKY130_FD_SC_HD__CLKBUF_1
XINPUT266 LA_IENA_MPRJ[105] VSSD VSSD VCCD VCCD NET266 SKY130_FD_SC_HD__CLKBUF_1
XINPUT267 LA_IENA_MPRJ[106] VSSD VSSD VCCD VCCD NET267 SKY130_FD_SC_HD__CLKBUF_1
XINPUT268 LA_IENA_MPRJ[107] VSSD VSSD VCCD VCCD NET268 SKY130_FD_SC_HD__CLKBUF_1
XINPUT269 LA_IENA_MPRJ[108] VSSD VSSD VCCD VCCD NET269 SKY130_FD_SC_HD__CLKBUF_1
XINPUT27 LA_DATA_OUT_CORE[120] VSSD VSSD VCCD VCCD NET27 SKY130_FD_SC_HD__BUF_2
XINPUT270 LA_IENA_MPRJ[109] VSSD VSSD VCCD VCCD NET270 SKY130_FD_SC_HD__CLKBUF_1
XINPUT271 LA_IENA_MPRJ[10] VSSD VSSD VCCD VCCD NET271 SKY130_FD_SC_HD__BUF_2
XINPUT272 LA_IENA_MPRJ[110] VSSD VSSD VCCD VCCD NET272 SKY130_FD_SC_HD__CLKBUF_1
XINPUT273 LA_IENA_MPRJ[111] VSSD VSSD VCCD VCCD NET273 SKY130_FD_SC_HD__CLKBUF_1
XINPUT274 LA_IENA_MPRJ[112] VSSD VSSD VCCD VCCD NET274 SKY130_FD_SC_HD__CLKBUF_1
XINPUT275 LA_IENA_MPRJ[113] VSSD VSSD VCCD VCCD NET275 SKY130_FD_SC_HD__CLKBUF_1
XINPUT276 LA_IENA_MPRJ[114] VSSD VSSD VCCD VCCD NET276 SKY130_FD_SC_HD__CLKBUF_1
XINPUT277 LA_IENA_MPRJ[115] VSSD VSSD VCCD VCCD NET277 SKY130_FD_SC_HD__CLKBUF_1
XINPUT278 LA_IENA_MPRJ[116] VSSD VSSD VCCD VCCD NET278 SKY130_FD_SC_HD__CLKBUF_1
XINPUT279 LA_IENA_MPRJ[117] VSSD VSSD VCCD VCCD NET279 SKY130_FD_SC_HD__CLKBUF_1
XINPUT28 LA_DATA_OUT_CORE[121] VSSD VSSD VCCD VCCD NET28 SKY130_FD_SC_HD__CLKBUF_4
XINPUT280 LA_IENA_MPRJ[118] VSSD VSSD VCCD VCCD NET280 SKY130_FD_SC_HD__CLKBUF_1
XINPUT281 LA_IENA_MPRJ[119] VSSD VSSD VCCD VCCD NET281 SKY130_FD_SC_HD__CLKBUF_1
XINPUT282 LA_IENA_MPRJ[11] VSSD VSSD VCCD VCCD NET282 SKY130_FD_SC_HD__CLKBUF_2
XINPUT283 LA_IENA_MPRJ[120] VSSD VSSD VCCD VCCD NET283 SKY130_FD_SC_HD__CLKBUF_1
XINPUT284 LA_IENA_MPRJ[121] VSSD VSSD VCCD VCCD NET284 SKY130_FD_SC_HD__CLKBUF_1
XINPUT285 LA_IENA_MPRJ[122] VSSD VSSD VCCD VCCD NET285 SKY130_FD_SC_HD__CLKBUF_1
XINPUT286 LA_IENA_MPRJ[123] VSSD VSSD VCCD VCCD NET286 SKY130_FD_SC_HD__CLKBUF_1
XINPUT287 LA_IENA_MPRJ[124] VSSD VSSD VCCD VCCD NET287 SKY130_FD_SC_HD__CLKBUF_1
XINPUT288 LA_IENA_MPRJ[125] VSSD VSSD VCCD VCCD NET288 SKY130_FD_SC_HD__CLKBUF_1
XINPUT289 LA_IENA_MPRJ[126] VSSD VSSD VCCD VCCD NET289 SKY130_FD_SC_HD__CLKBUF_1
XINPUT29 LA_DATA_OUT_CORE[122] VSSD VSSD VCCD VCCD NET29 SKY130_FD_SC_HD__BUF_4
XINPUT290 LA_IENA_MPRJ[127] VSSD VSSD VCCD VCCD NET290 SKY130_FD_SC_HD__CLKBUF_1
XINPUT291 LA_IENA_MPRJ[12] VSSD VSSD VCCD VCCD NET291 SKY130_FD_SC_HD__BUF_2
XINPUT292 LA_IENA_MPRJ[13] VSSD VSSD VCCD VCCD NET292 SKY130_FD_SC_HD__CLKBUF_1
XINPUT293 LA_IENA_MPRJ[14] VSSD VSSD VCCD VCCD NET293 SKY130_FD_SC_HD__CLKBUF_1
XINPUT294 LA_IENA_MPRJ[15] VSSD VSSD VCCD VCCD NET294 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT295 LA_IENA_MPRJ[16] VSSD VSSD VCCD VCCD NET295 SKY130_FD_SC_HD__CLKBUF_1
XINPUT296 LA_IENA_MPRJ[17] VSSD VSSD VCCD VCCD NET296 SKY130_FD_SC_HD__CLKBUF_1
XINPUT297 LA_IENA_MPRJ[18] VSSD VSSD VCCD VCCD NET297 SKY130_FD_SC_HD__CLKBUF_1
XINPUT298 LA_IENA_MPRJ[19] VSSD VSSD VCCD VCCD NET298 SKY130_FD_SC_HD__CLKBUF_1
XINPUT299 LA_IENA_MPRJ[1] VSSD VSSD VCCD VCCD NET299 SKY130_FD_SC_HD__CLKBUF_1
XINPUT3 CARAVEL_RSTN VSSD VSSD VCCD VCCD NET3 SKY130_FD_SC_HD__CLKBUF_1
XINPUT30 LA_DATA_OUT_CORE[123] VSSD VSSD VCCD VCCD NET30 SKY130_FD_SC_HD__CLKBUF_4
XINPUT300 LA_IENA_MPRJ[20] VSSD VSSD VCCD VCCD NET300 SKY130_FD_SC_HD__CLKBUF_1
XINPUT301 LA_IENA_MPRJ[21] VSSD VSSD VCCD VCCD NET301 SKY130_FD_SC_HD__CLKBUF_1
XINPUT302 LA_IENA_MPRJ[22] VSSD VSSD VCCD VCCD NET302 SKY130_FD_SC_HD__CLKBUF_1
XINPUT303 LA_IENA_MPRJ[23] VSSD VSSD VCCD VCCD NET303 SKY130_FD_SC_HD__CLKBUF_1
XINPUT304 LA_IENA_MPRJ[24] VSSD VSSD VCCD VCCD NET304 SKY130_FD_SC_HD__CLKBUF_1
XINPUT305 LA_IENA_MPRJ[25] VSSD VSSD VCCD VCCD NET305 SKY130_FD_SC_HD__CLKBUF_1
XINPUT306 LA_IENA_MPRJ[26] VSSD VSSD VCCD VCCD NET306 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT307 LA_IENA_MPRJ[27] VSSD VSSD VCCD VCCD NET307 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT308 LA_IENA_MPRJ[28] VSSD VSSD VCCD VCCD NET308 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT309 LA_IENA_MPRJ[29] VSSD VSSD VCCD VCCD NET309 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT31 LA_DATA_OUT_CORE[124] VSSD VSSD VCCD VCCD NET31 SKY130_FD_SC_HD__CLKBUF_4
XINPUT310 LA_IENA_MPRJ[2] VSSD VSSD VCCD VCCD NET310 SKY130_FD_SC_HD__CLKBUF_1
XINPUT311 LA_IENA_MPRJ[30] VSSD VSSD VCCD VCCD NET311 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT312 LA_IENA_MPRJ[31] VSSD VSSD VCCD VCCD NET312 SKY130_FD_SC_HD__CLKBUF_1
XINPUT313 LA_IENA_MPRJ[32] VSSD VSSD VCCD VCCD NET313 SKY130_FD_SC_HD__CLKBUF_1
XINPUT314 LA_IENA_MPRJ[33] VSSD VSSD VCCD VCCD NET314 SKY130_FD_SC_HD__CLKBUF_1
XINPUT315 LA_IENA_MPRJ[34] VSSD VSSD VCCD VCCD NET315 SKY130_FD_SC_HD__CLKBUF_1
XINPUT316 LA_IENA_MPRJ[35] VSSD VSSD VCCD VCCD NET316 SKY130_FD_SC_HD__CLKBUF_1
XINPUT317 LA_IENA_MPRJ[36] VSSD VSSD VCCD VCCD NET317 SKY130_FD_SC_HD__CLKBUF_1
XINPUT318 LA_IENA_MPRJ[37] VSSD VSSD VCCD VCCD NET318 SKY130_FD_SC_HD__CLKBUF_1
XINPUT319 LA_IENA_MPRJ[38] VSSD VSSD VCCD VCCD NET319 SKY130_FD_SC_HD__CLKBUF_1
XINPUT32 LA_DATA_OUT_CORE[125] VSSD VSSD VCCD VCCD NET32 SKY130_FD_SC_HD__CLKBUF_4
XINPUT320 LA_IENA_MPRJ[39] VSSD VSSD VCCD VCCD NET320 SKY130_FD_SC_HD__CLKBUF_1
XINPUT321 LA_IENA_MPRJ[3] VSSD VSSD VCCD VCCD NET321 SKY130_FD_SC_HD__CLKBUF_1
XINPUT322 LA_IENA_MPRJ[40] VSSD VSSD VCCD VCCD NET322 SKY130_FD_SC_HD__CLKBUF_1
XINPUT323 LA_IENA_MPRJ[41] VSSD VSSD VCCD VCCD NET323 SKY130_FD_SC_HD__CLKBUF_1
XINPUT324 LA_IENA_MPRJ[42] VSSD VSSD VCCD VCCD NET324 SKY130_FD_SC_HD__CLKBUF_1
XINPUT325 LA_IENA_MPRJ[43] VSSD VSSD VCCD VCCD NET325 SKY130_FD_SC_HD__CLKBUF_1
XINPUT326 LA_IENA_MPRJ[44] VSSD VSSD VCCD VCCD NET326 SKY130_FD_SC_HD__CLKBUF_1
XINPUT327 LA_IENA_MPRJ[45] VSSD VSSD VCCD VCCD NET327 SKY130_FD_SC_HD__CLKBUF_1
XINPUT328 LA_IENA_MPRJ[46] VSSD VSSD VCCD VCCD NET328 SKY130_FD_SC_HD__CLKBUF_1
XINPUT329 LA_IENA_MPRJ[47] VSSD VSSD VCCD VCCD NET329 SKY130_FD_SC_HD__CLKBUF_1
XINPUT33 LA_DATA_OUT_CORE[126] VSSD VSSD VCCD VCCD NET33 SKY130_FD_SC_HD__CLKBUF_4
XINPUT330 LA_IENA_MPRJ[48] VSSD VSSD VCCD VCCD NET330 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT331 LA_IENA_MPRJ[49] VSSD VSSD VCCD VCCD NET331 SKY130_FD_SC_HD__CLKBUF_1
XINPUT332 LA_IENA_MPRJ[4] VSSD VSSD VCCD VCCD NET332 SKY130_FD_SC_HD__CLKBUF_1
XINPUT333 LA_IENA_MPRJ[50] VSSD VSSD VCCD VCCD NET333 SKY130_FD_SC_HD__CLKBUF_1
XINPUT334 LA_IENA_MPRJ[51] VSSD VSSD VCCD VCCD NET334 SKY130_FD_SC_HD__CLKBUF_1
XINPUT335 LA_IENA_MPRJ[52] VSSD VSSD VCCD VCCD NET335 SKY130_FD_SC_HD__CLKBUF_1
XINPUT336 LA_IENA_MPRJ[53] VSSD VSSD VCCD VCCD NET336 SKY130_FD_SC_HD__CLKBUF_1
XINPUT337 LA_IENA_MPRJ[54] VSSD VSSD VCCD VCCD NET337 SKY130_FD_SC_HD__CLKBUF_1
XINPUT338 LA_IENA_MPRJ[55] VSSD VSSD VCCD VCCD NET338 SKY130_FD_SC_HD__CLKBUF_1
XINPUT339 LA_IENA_MPRJ[56] VSSD VSSD VCCD VCCD NET339 SKY130_FD_SC_HD__CLKBUF_1
XINPUT34 LA_DATA_OUT_CORE[127] VSSD VSSD VCCD VCCD NET34 SKY130_FD_SC_HD__CLKBUF_4
XINPUT340 LA_IENA_MPRJ[57] VSSD VSSD VCCD VCCD NET340 SKY130_FD_SC_HD__CLKBUF_1
XINPUT341 LA_IENA_MPRJ[58] VSSD VSSD VCCD VCCD NET341 SKY130_FD_SC_HD__CLKBUF_1
XINPUT342 LA_IENA_MPRJ[59] VSSD VSSD VCCD VCCD NET342 SKY130_FD_SC_HD__CLKBUF_1
XINPUT343 LA_IENA_MPRJ[5] VSSD VSSD VCCD VCCD NET343 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT344 LA_IENA_MPRJ[60] VSSD VSSD VCCD VCCD NET344 SKY130_FD_SC_HD__CLKBUF_1
XINPUT345 LA_IENA_MPRJ[61] VSSD VSSD VCCD VCCD NET345 SKY130_FD_SC_HD__CLKBUF_1
XINPUT346 LA_IENA_MPRJ[62] VSSD VSSD VCCD VCCD NET346 SKY130_FD_SC_HD__CLKBUF_1
XINPUT347 LA_IENA_MPRJ[63] VSSD VSSD VCCD VCCD NET347 SKY130_FD_SC_HD__CLKBUF_1
XINPUT348 LA_IENA_MPRJ[64] VSSD VSSD VCCD VCCD NET348 SKY130_FD_SC_HD__CLKBUF_1
XINPUT349 LA_IENA_MPRJ[65] VSSD VSSD VCCD VCCD NET349 SKY130_FD_SC_HD__CLKBUF_1
XINPUT35 LA_DATA_OUT_CORE[12] VSSD VSSD VCCD VCCD NET35 SKY130_FD_SC_HD__BUF_2
XINPUT350 LA_IENA_MPRJ[66] VSSD VSSD VCCD VCCD NET350 SKY130_FD_SC_HD__CLKBUF_1
XINPUT351 LA_IENA_MPRJ[67] VSSD VSSD VCCD VCCD NET351 SKY130_FD_SC_HD__CLKBUF_1
XINPUT352 LA_IENA_MPRJ[68] VSSD VSSD VCCD VCCD NET352 SKY130_FD_SC_HD__CLKBUF_1
XINPUT353 LA_IENA_MPRJ[69] VSSD VSSD VCCD VCCD NET353 SKY130_FD_SC_HD__CLKBUF_1
XINPUT354 LA_IENA_MPRJ[6] VSSD VSSD VCCD VCCD NET354 SKY130_FD_SC_HD__CLKBUF_1
XINPUT355 LA_IENA_MPRJ[70] VSSD VSSD VCCD VCCD NET355 SKY130_FD_SC_HD__CLKBUF_1
XINPUT356 LA_IENA_MPRJ[71] VSSD VSSD VCCD VCCD NET356 SKY130_FD_SC_HD__CLKBUF_1
XINPUT357 LA_IENA_MPRJ[72] VSSD VSSD VCCD VCCD NET357 SKY130_FD_SC_HD__CLKBUF_1
XINPUT358 LA_IENA_MPRJ[73] VSSD VSSD VCCD VCCD NET358 SKY130_FD_SC_HD__CLKBUF_1
XINPUT359 LA_IENA_MPRJ[74] VSSD VSSD VCCD VCCD NET359 SKY130_FD_SC_HD__CLKBUF_1
XINPUT36 LA_DATA_OUT_CORE[13] VSSD VSSD VCCD VCCD NET36 SKY130_FD_SC_HD__CLKBUF_4
XINPUT360 LA_IENA_MPRJ[75] VSSD VSSD VCCD VCCD NET360 SKY130_FD_SC_HD__CLKBUF_1
XINPUT361 LA_IENA_MPRJ[76] VSSD VSSD VCCD VCCD NET361 SKY130_FD_SC_HD__CLKBUF_1
XINPUT362 LA_IENA_MPRJ[77] VSSD VSSD VCCD VCCD NET362 SKY130_FD_SC_HD__CLKBUF_1
XINPUT363 LA_IENA_MPRJ[78] VSSD VSSD VCCD VCCD NET363 SKY130_FD_SC_HD__CLKBUF_1
XINPUT364 LA_IENA_MPRJ[79] VSSD VSSD VCCD VCCD NET364 SKY130_FD_SC_HD__CLKBUF_1
XINPUT365 LA_IENA_MPRJ[7] VSSD VSSD VCCD VCCD NET365 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT366 LA_IENA_MPRJ[80] VSSD VSSD VCCD VCCD NET366 SKY130_FD_SC_HD__CLKBUF_1
XINPUT367 LA_IENA_MPRJ[81] VSSD VSSD VCCD VCCD NET367 SKY130_FD_SC_HD__CLKBUF_1
XINPUT368 LA_IENA_MPRJ[82] VSSD VSSD VCCD VCCD NET368 SKY130_FD_SC_HD__CLKBUF_1
XINPUT369 LA_IENA_MPRJ[83] VSSD VSSD VCCD VCCD NET369 SKY130_FD_SC_HD__CLKBUF_1
XINPUT37 LA_DATA_OUT_CORE[14] VSSD VSSD VCCD VCCD NET37 SKY130_FD_SC_HD__BUF_4
XINPUT370 LA_IENA_MPRJ[84] VSSD VSSD VCCD VCCD NET370 SKY130_FD_SC_HD__CLKBUF_1
XINPUT371 LA_IENA_MPRJ[85] VSSD VSSD VCCD VCCD NET371 SKY130_FD_SC_HD__CLKBUF_1
XINPUT372 LA_IENA_MPRJ[86] VSSD VSSD VCCD VCCD NET372 SKY130_FD_SC_HD__CLKBUF_1
XINPUT373 LA_IENA_MPRJ[87] VSSD VSSD VCCD VCCD NET373 SKY130_FD_SC_HD__CLKBUF_1
XINPUT374 LA_IENA_MPRJ[88] VSSD VSSD VCCD VCCD NET374 SKY130_FD_SC_HD__CLKBUF_1
XINPUT375 LA_IENA_MPRJ[89] VSSD VSSD VCCD VCCD NET375 SKY130_FD_SC_HD__CLKBUF_1
XINPUT376 LA_IENA_MPRJ[8] VSSD VSSD VCCD VCCD NET376 SKY130_FD_SC_HD__CLKBUF_2
XINPUT377 LA_IENA_MPRJ[90] VSSD VSSD VCCD VCCD NET377 SKY130_FD_SC_HD__CLKBUF_1
XINPUT378 LA_IENA_MPRJ[91] VSSD VSSD VCCD VCCD NET378 SKY130_FD_SC_HD__CLKBUF_1
XINPUT379 LA_IENA_MPRJ[92] VSSD VSSD VCCD VCCD NET379 SKY130_FD_SC_HD__CLKBUF_1
XINPUT38 LA_DATA_OUT_CORE[15] VSSD VSSD VCCD VCCD NET38 SKY130_FD_SC_HD__BUF_4
XINPUT380 LA_IENA_MPRJ[93] VSSD VSSD VCCD VCCD NET380 SKY130_FD_SC_HD__CLKBUF_1
XINPUT381 LA_IENA_MPRJ[94] VSSD VSSD VCCD VCCD NET381 SKY130_FD_SC_HD__CLKBUF_1
XINPUT382 LA_IENA_MPRJ[95] VSSD VSSD VCCD VCCD NET382 SKY130_FD_SC_HD__CLKBUF_1
XINPUT383 LA_IENA_MPRJ[96] VSSD VSSD VCCD VCCD NET383 SKY130_FD_SC_HD__CLKBUF_1
XINPUT384 LA_IENA_MPRJ[97] VSSD VSSD VCCD VCCD NET384 SKY130_FD_SC_HD__CLKBUF_1
XINPUT385 LA_IENA_MPRJ[98] VSSD VSSD VCCD VCCD NET385 SKY130_FD_SC_HD__CLKBUF_1
XINPUT386 LA_IENA_MPRJ[99] VSSD VSSD VCCD VCCD NET386 SKY130_FD_SC_HD__CLKBUF_1
XINPUT387 LA_IENA_MPRJ[9] VSSD VSSD VCCD VCCD NET387 SKY130_FD_SC_HD__CLKBUF_2
XINPUT388 LA_OENB_MPRJ[0] VSSD VSSD VCCD VCCD NET388 SKY130_FD_SC_HD__CLKBUF_2
XINPUT389 LA_OENB_MPRJ[100] VSSD VSSD VCCD VCCD NET389 SKY130_FD_SC_HD__CLKBUF_4
XINPUT39 LA_DATA_OUT_CORE[16] VSSD VSSD VCCD VCCD NET39 SKY130_FD_SC_HD__BUF_4
XINPUT390 LA_OENB_MPRJ[101] VSSD VSSD VCCD VCCD NET390 SKY130_FD_SC_HD__CLKBUF_4
XINPUT391 LA_OENB_MPRJ[102] VSSD VSSD VCCD VCCD NET391 SKY130_FD_SC_HD__CLKBUF_4
XINPUT392 LA_OENB_MPRJ[103] VSSD VSSD VCCD VCCD NET392 SKY130_FD_SC_HD__CLKBUF_4
XINPUT393 LA_OENB_MPRJ[104] VSSD VSSD VCCD VCCD NET393 SKY130_FD_SC_HD__CLKBUF_2
XINPUT394 LA_OENB_MPRJ[105] VSSD VSSD VCCD VCCD NET394 SKY130_FD_SC_HD__BUF_2
XINPUT395 LA_OENB_MPRJ[106] VSSD VSSD VCCD VCCD NET395 SKY130_FD_SC_HD__CLKBUF_4
XINPUT396 LA_OENB_MPRJ[107] VSSD VSSD VCCD VCCD NET396 SKY130_FD_SC_HD__CLKBUF_4
XINPUT397 LA_OENB_MPRJ[108] VSSD VSSD VCCD VCCD NET397 SKY130_FD_SC_HD__BUF_2
XINPUT398 LA_OENB_MPRJ[109] VSSD VSSD VCCD VCCD NET398 SKY130_FD_SC_HD__CLKBUF_4
XINPUT399 LA_OENB_MPRJ[10] VSSD VSSD VCCD VCCD NET399 SKY130_FD_SC_HD__CLKBUF_2
XINPUT4 LA_DATA_OUT_CORE[0] VSSD VSSD VCCD VCCD NET4 SKY130_FD_SC_HD__BUF_4
XINPUT40 LA_DATA_OUT_CORE[17] VSSD VSSD VCCD VCCD NET40 SKY130_FD_SC_HD__CLKBUF_4
XINPUT400 LA_OENB_MPRJ[110] VSSD VSSD VCCD VCCD NET400 SKY130_FD_SC_HD__CLKBUF_4
XINPUT401 LA_OENB_MPRJ[111] VSSD VSSD VCCD VCCD NET401 SKY130_FD_SC_HD__CLKBUF_4
XINPUT402 LA_OENB_MPRJ[112] VSSD VSSD VCCD VCCD NET402 SKY130_FD_SC_HD__BUF_2
XINPUT403 LA_OENB_MPRJ[113] VSSD VSSD VCCD VCCD NET403 SKY130_FD_SC_HD__CLKBUF_4
XINPUT404 LA_OENB_MPRJ[114] VSSD VSSD VCCD VCCD NET404 SKY130_FD_SC_HD__CLKBUF_4
XINPUT405 LA_OENB_MPRJ[115] VSSD VSSD VCCD VCCD NET405 SKY130_FD_SC_HD__CLKBUF_4
XINPUT406 LA_OENB_MPRJ[116] VSSD VSSD VCCD VCCD NET406 SKY130_FD_SC_HD__CLKBUF_4
XINPUT407 LA_OENB_MPRJ[117] VSSD VSSD VCCD VCCD NET407 SKY130_FD_SC_HD__CLKBUF_4
XINPUT408 LA_OENB_MPRJ[118] VSSD VSSD VCCD VCCD NET408 SKY130_FD_SC_HD__CLKBUF_4
XINPUT409 LA_OENB_MPRJ[119] VSSD VSSD VCCD VCCD NET409 SKY130_FD_SC_HD__CLKBUF_4
XINPUT41 LA_DATA_OUT_CORE[18] VSSD VSSD VCCD VCCD NET41 SKY130_FD_SC_HD__CLKBUF_4
XINPUT410 LA_OENB_MPRJ[11] VSSD VSSD VCCD VCCD NET410 SKY130_FD_SC_HD__CLKBUF_2
XINPUT411 LA_OENB_MPRJ[120] VSSD VSSD VCCD VCCD NET411 SKY130_FD_SC_HD__CLKBUF_4
XINPUT412 LA_OENB_MPRJ[121] VSSD VSSD VCCD VCCD NET412 SKY130_FD_SC_HD__BUF_2
XINPUT413 LA_OENB_MPRJ[122] VSSD VSSD VCCD VCCD NET413 SKY130_FD_SC_HD__BUF_2
XINPUT414 LA_OENB_MPRJ[123] VSSD VSSD VCCD VCCD NET414 SKY130_FD_SC_HD__CLKBUF_4
XINPUT415 LA_OENB_MPRJ[124] VSSD VSSD VCCD VCCD NET415 SKY130_FD_SC_HD__CLKBUF_4
XINPUT416 LA_OENB_MPRJ[125] VSSD VSSD VCCD VCCD NET416 SKY130_FD_SC_HD__CLKBUF_4
XINPUT417 LA_OENB_MPRJ[126] VSSD VSSD VCCD VCCD NET417 SKY130_FD_SC_HD__CLKBUF_4
XINPUT418 LA_OENB_MPRJ[127] VSSD VSSD VCCD VCCD NET418 SKY130_FD_SC_HD__BUF_2
XINPUT419 LA_OENB_MPRJ[12] VSSD VSSD VCCD VCCD NET419 SKY130_FD_SC_HD__CLKBUF_2
XINPUT42 LA_DATA_OUT_CORE[19] VSSD VSSD VCCD VCCD NET42 SKY130_FD_SC_HD__CLKBUF_4
XINPUT420 LA_OENB_MPRJ[13] VSSD VSSD VCCD VCCD NET420 SKY130_FD_SC_HD__BUF_2
XINPUT421 LA_OENB_MPRJ[14] VSSD VSSD VCCD VCCD NET421 SKY130_FD_SC_HD__CLKBUF_4
XINPUT422 LA_OENB_MPRJ[15] VSSD VSSD VCCD VCCD NET422 SKY130_FD_SC_HD__BUF_2
XINPUT423 LA_OENB_MPRJ[16] VSSD VSSD VCCD VCCD NET423 SKY130_FD_SC_HD__CLKBUF_2
XINPUT424 LA_OENB_MPRJ[17] VSSD VSSD VCCD VCCD NET424 SKY130_FD_SC_HD__BUF_2
XINPUT425 LA_OENB_MPRJ[18] VSSD VSSD VCCD VCCD NET425 SKY130_FD_SC_HD__CLKBUF_2
XINPUT426 LA_OENB_MPRJ[19] VSSD VSSD VCCD VCCD NET426 SKY130_FD_SC_HD__CLKBUF_4
XINPUT427 LA_OENB_MPRJ[1] VSSD VSSD VCCD VCCD NET427 SKY130_FD_SC_HD__CLKBUF_2
XINPUT428 LA_OENB_MPRJ[20] VSSD VSSD VCCD VCCD NET428 SKY130_FD_SC_HD__CLKBUF_4
XINPUT429 LA_OENB_MPRJ[21] VSSD VSSD VCCD VCCD NET429 SKY130_FD_SC_HD__BUF_2
XINPUT43 LA_DATA_OUT_CORE[1] VSSD VSSD VCCD VCCD NET43 SKY130_FD_SC_HD__BUF_4
XINPUT430 LA_OENB_MPRJ[22] VSSD VSSD VCCD VCCD NET430 SKY130_FD_SC_HD__CLKBUF_4
XINPUT431 LA_OENB_MPRJ[23] VSSD VSSD VCCD VCCD NET431 SKY130_FD_SC_HD__BUF_2
XINPUT432 LA_OENB_MPRJ[24] VSSD VSSD VCCD VCCD NET432 SKY130_FD_SC_HD__BUF_2
XINPUT433 LA_OENB_MPRJ[25] VSSD VSSD VCCD VCCD NET433 SKY130_FD_SC_HD__BUF_2
XINPUT434 LA_OENB_MPRJ[26] VSSD VSSD VCCD VCCD NET434 SKY130_FD_SC_HD__BUF_2
XINPUT435 LA_OENB_MPRJ[27] VSSD VSSD VCCD VCCD NET435 SKY130_FD_SC_HD__BUF_2
XINPUT436 LA_OENB_MPRJ[28] VSSD VSSD VCCD VCCD NET436 SKY130_FD_SC_HD__BUF_2
XINPUT437 LA_OENB_MPRJ[29] VSSD VSSD VCCD VCCD NET437 SKY130_FD_SC_HD__BUF_2
XINPUT438 LA_OENB_MPRJ[2] VSSD VSSD VCCD VCCD NET438 SKY130_FD_SC_HD__BUF_2
XINPUT439 LA_OENB_MPRJ[30] VSSD VSSD VCCD VCCD NET439 SKY130_FD_SC_HD__CLKBUF_2
XINPUT44 LA_DATA_OUT_CORE[20] VSSD VSSD VCCD VCCD NET44 SKY130_FD_SC_HD__CLKBUF_4
XINPUT440 LA_OENB_MPRJ[31] VSSD VSSD VCCD VCCD NET440 SKY130_FD_SC_HD__BUF_2
XINPUT441 LA_OENB_MPRJ[32] VSSD VSSD VCCD VCCD NET441 SKY130_FD_SC_HD__BUF_2
XINPUT442 LA_OENB_MPRJ[33] VSSD VSSD VCCD VCCD NET442 SKY130_FD_SC_HD__BUF_2
XINPUT443 LA_OENB_MPRJ[34] VSSD VSSD VCCD VCCD NET443 SKY130_FD_SC_HD__CLKBUF_2
XINPUT444 LA_OENB_MPRJ[35] VSSD VSSD VCCD VCCD NET444 SKY130_FD_SC_HD__CLKBUF_2
XINPUT445 LA_OENB_MPRJ[36] VSSD VSSD VCCD VCCD NET445 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT446 LA_OENB_MPRJ[37] VSSD VSSD VCCD VCCD NET446 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT447 LA_OENB_MPRJ[38] VSSD VSSD VCCD VCCD NET447 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT448 LA_OENB_MPRJ[39] VSSD VSSD VCCD VCCD NET448 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT449 LA_OENB_MPRJ[3] VSSD VSSD VCCD VCCD NET449 SKY130_FD_SC_HD__CLKBUF_2
XINPUT45 LA_DATA_OUT_CORE[21] VSSD VSSD VCCD VCCD NET45 SKY130_FD_SC_HD__CLKBUF_4
XINPUT450 LA_OENB_MPRJ[40] VSSD VSSD VCCD VCCD NET450 SKY130_FD_SC_HD__BUF_4
XINPUT451 LA_OENB_MPRJ[41] VSSD VSSD VCCD VCCD NET451 SKY130_FD_SC_HD__CLKBUF_2
XINPUT452 LA_OENB_MPRJ[42] VSSD VSSD VCCD VCCD NET452 SKY130_FD_SC_HD__BUF_4
XINPUT453 LA_OENB_MPRJ[43] VSSD VSSD VCCD VCCD NET453 SKY130_FD_SC_HD__BUF_4
XINPUT454 LA_OENB_MPRJ[44] VSSD VSSD VCCD VCCD NET454 SKY130_FD_SC_HD__CLKBUF_2
XINPUT455 LA_OENB_MPRJ[45] VSSD VSSD VCCD VCCD NET455 SKY130_FD_SC_HD__CLKBUF_2
XINPUT456 LA_OENB_MPRJ[46] VSSD VSSD VCCD VCCD NET456 SKY130_FD_SC_HD__CLKBUF_2
XINPUT457 LA_OENB_MPRJ[47] VSSD VSSD VCCD VCCD NET457 SKY130_FD_SC_HD__BUF_4
XINPUT458 LA_OENB_MPRJ[48] VSSD VSSD VCCD VCCD NET458 SKY130_FD_SC_HD__CLKBUF_2
XINPUT459 LA_OENB_MPRJ[49] VSSD VSSD VCCD VCCD NET459 SKY130_FD_SC_HD__BUF_2
XINPUT46 LA_DATA_OUT_CORE[22] VSSD VSSD VCCD VCCD NET46 SKY130_FD_SC_HD__CLKBUF_4
XINPUT460 LA_OENB_MPRJ[4] VSSD VSSD VCCD VCCD NET460 SKY130_FD_SC_HD__CLKBUF_2
XINPUT461 LA_OENB_MPRJ[50] VSSD VSSD VCCD VCCD NET461 SKY130_FD_SC_HD__CLKBUF_2
XINPUT462 LA_OENB_MPRJ[51] VSSD VSSD VCCD VCCD NET462 SKY130_FD_SC_HD__CLKBUF_2
XINPUT463 LA_OENB_MPRJ[52] VSSD VSSD VCCD VCCD NET463 SKY130_FD_SC_HD__CLKBUF_2
XINPUT464 LA_OENB_MPRJ[53] VSSD VSSD VCCD VCCD NET464 SKY130_FD_SC_HD__BUF_2
XINPUT465 LA_OENB_MPRJ[54] VSSD VSSD VCCD VCCD NET465 SKY130_FD_SC_HD__CLKBUF_2
XINPUT466 LA_OENB_MPRJ[55] VSSD VSSD VCCD VCCD NET466 SKY130_FD_SC_HD__BUF_2
XINPUT467 LA_OENB_MPRJ[56] VSSD VSSD VCCD VCCD NET467 SKY130_FD_SC_HD__CLKBUF_2
XINPUT468 LA_OENB_MPRJ[57] VSSD VSSD VCCD VCCD NET468 SKY130_FD_SC_HD__BUF_2
XINPUT469 LA_OENB_MPRJ[58] VSSD VSSD VCCD VCCD NET469 SKY130_FD_SC_HD__CLKBUF_2
XINPUT47 LA_DATA_OUT_CORE[23] VSSD VSSD VCCD VCCD NET47 SKY130_FD_SC_HD__CLKBUF_4
XINPUT470 LA_OENB_MPRJ[59] VSSD VSSD VCCD VCCD NET470 SKY130_FD_SC_HD__BUF_2
XINPUT471 LA_OENB_MPRJ[5] VSSD VSSD VCCD VCCD NET471 SKY130_FD_SC_HD__CLKBUF_2
XINPUT472 LA_OENB_MPRJ[60] VSSD VSSD VCCD VCCD NET472 SKY130_FD_SC_HD__CLKBUF_2
XINPUT473 LA_OENB_MPRJ[61] VSSD VSSD VCCD VCCD NET473 SKY130_FD_SC_HD__CLKBUF_2
XINPUT474 LA_OENB_MPRJ[62] VSSD VSSD VCCD VCCD NET474 SKY130_FD_SC_HD__CLKBUF_2
XINPUT475 LA_OENB_MPRJ[63] VSSD VSSD VCCD VCCD NET475 SKY130_FD_SC_HD__BUF_2
XINPUT476 LA_OENB_MPRJ[64] VSSD VSSD VCCD VCCD NET476 SKY130_FD_SC_HD__BUF_2
XINPUT477 LA_OENB_MPRJ[65] VSSD VSSD VCCD VCCD NET477 SKY130_FD_SC_HD__BUF_2
XINPUT478 LA_OENB_MPRJ[66] VSSD VSSD VCCD VCCD NET478 SKY130_FD_SC_HD__BUF_4
XINPUT479 LA_OENB_MPRJ[67] VSSD VSSD VCCD VCCD NET479 SKY130_FD_SC_HD__BUF_2
XINPUT48 LA_DATA_OUT_CORE[24] VSSD VSSD VCCD VCCD NET48 SKY130_FD_SC_HD__CLKBUF_4
XINPUT480 LA_OENB_MPRJ[68] VSSD VSSD VCCD VCCD NET480 SKY130_FD_SC_HD__CLKBUF_2
XINPUT481 LA_OENB_MPRJ[69] VSSD VSSD VCCD VCCD NET481 SKY130_FD_SC_HD__BUF_2
XINPUT482 LA_OENB_MPRJ[6] VSSD VSSD VCCD VCCD NET482 SKY130_FD_SC_HD__CLKBUF_2
XINPUT483 LA_OENB_MPRJ[70] VSSD VSSD VCCD VCCD NET483 SKY130_FD_SC_HD__BUF_2
XINPUT484 LA_OENB_MPRJ[71] VSSD VSSD VCCD VCCD NET484 SKY130_FD_SC_HD__CLKBUF_2
XINPUT485 LA_OENB_MPRJ[72] VSSD VSSD VCCD VCCD NET485 SKY130_FD_SC_HD__BUF_2
XINPUT486 LA_OENB_MPRJ[73] VSSD VSSD VCCD VCCD NET486 SKY130_FD_SC_HD__BUF_2
XINPUT487 LA_OENB_MPRJ[74] VSSD VSSD VCCD VCCD NET487 SKY130_FD_SC_HD__BUF_2
XINPUT488 LA_OENB_MPRJ[75] VSSD VSSD VCCD VCCD NET488 SKY130_FD_SC_HD__BUF_2
XINPUT489 LA_OENB_MPRJ[76] VSSD VSSD VCCD VCCD NET489 SKY130_FD_SC_HD__CLKBUF_4
XINPUT49 LA_DATA_OUT_CORE[25] VSSD VSSD VCCD VCCD NET49 SKY130_FD_SC_HD__CLKBUF_4
XINPUT490 LA_OENB_MPRJ[77] VSSD VSSD VCCD VCCD NET490 SKY130_FD_SC_HD__BUF_2
XINPUT491 LA_OENB_MPRJ[78] VSSD VSSD VCCD VCCD NET491 SKY130_FD_SC_HD__CLKBUF_4
XINPUT492 LA_OENB_MPRJ[79] VSSD VSSD VCCD VCCD NET492 SKY130_FD_SC_HD__CLKBUF_4
XINPUT493 LA_OENB_MPRJ[7] VSSD VSSD VCCD VCCD NET493 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT494 LA_OENB_MPRJ[80] VSSD VSSD VCCD VCCD NET494 SKY130_FD_SC_HD__BUF_4
XINPUT495 LA_OENB_MPRJ[81] VSSD VSSD VCCD VCCD NET495 SKY130_FD_SC_HD__CLKBUF_4
XINPUT496 LA_OENB_MPRJ[82] VSSD VSSD VCCD VCCD NET496 SKY130_FD_SC_HD__BUF_4
XINPUT497 LA_OENB_MPRJ[83] VSSD VSSD VCCD VCCD NET497 SKY130_FD_SC_HD__BUF_4
XINPUT498 LA_OENB_MPRJ[84] VSSD VSSD VCCD VCCD NET498 SKY130_FD_SC_HD__BUF_4
XINPUT499 LA_OENB_MPRJ[85] VSSD VSSD VCCD VCCD NET499 SKY130_FD_SC_HD__BUF_4
XINPUT5 LA_DATA_OUT_CORE[100] VSSD VSSD VCCD VCCD NET5 SKY130_FD_SC_HD__BUF_4
XINPUT50 LA_DATA_OUT_CORE[26] VSSD VSSD VCCD VCCD NET50 SKY130_FD_SC_HD__CLKBUF_4
XINPUT500 LA_OENB_MPRJ[86] VSSD VSSD VCCD VCCD NET500 SKY130_FD_SC_HD__CLKBUF_4
XINPUT501 LA_OENB_MPRJ[87] VSSD VSSD VCCD VCCD NET501 SKY130_FD_SC_HD__CLKBUF_4
XINPUT502 LA_OENB_MPRJ[88] VSSD VSSD VCCD VCCD NET502 SKY130_FD_SC_HD__CLKBUF_4
XINPUT503 LA_OENB_MPRJ[89] VSSD VSSD VCCD VCCD NET503 SKY130_FD_SC_HD__CLKBUF_4
XINPUT504 LA_OENB_MPRJ[8] VSSD VSSD VCCD VCCD NET504 SKY130_FD_SC_HD__BUF_2
XINPUT505 LA_OENB_MPRJ[90] VSSD VSSD VCCD VCCD NET505 SKY130_FD_SC_HD__BUF_2
XINPUT506 LA_OENB_MPRJ[91] VSSD VSSD VCCD VCCD NET506 SKY130_FD_SC_HD__CLKBUF_4
XINPUT507 LA_OENB_MPRJ[92] VSSD VSSD VCCD VCCD NET507 SKY130_FD_SC_HD__BUF_2
XINPUT508 LA_OENB_MPRJ[93] VSSD VSSD VCCD VCCD NET508 SKY130_FD_SC_HD__BUF_2
XINPUT509 LA_OENB_MPRJ[94] VSSD VSSD VCCD VCCD NET509 SKY130_FD_SC_HD__BUF_2
XINPUT51 LA_DATA_OUT_CORE[27] VSSD VSSD VCCD VCCD NET51 SKY130_FD_SC_HD__CLKBUF_4
XINPUT510 LA_OENB_MPRJ[95] VSSD VSSD VCCD VCCD NET510 SKY130_FD_SC_HD__CLKBUF_4
XINPUT511 LA_OENB_MPRJ[96] VSSD VSSD VCCD VCCD NET511 SKY130_FD_SC_HD__CLKBUF_4
XINPUT512 LA_OENB_MPRJ[97] VSSD VSSD VCCD VCCD NET512 SKY130_FD_SC_HD__CLKBUF_4
XINPUT513 LA_OENB_MPRJ[98] VSSD VSSD VCCD VCCD NET513 SKY130_FD_SC_HD__CLKBUF_2
XINPUT514 LA_OENB_MPRJ[99] VSSD VSSD VCCD VCCD NET514 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT515 LA_OENB_MPRJ[9] VSSD VSSD VCCD VCCD NET515 SKY130_FD_SC_HD__CLKBUF_2
XINPUT516 MPRJ_ACK_I_USER VSSD VSSD VCCD VCCD NET516 SKY130_FD_SC_HD__BUF_12
XINPUT517 MPRJ_ADR_O_CORE[0] VSSD VSSD VCCD VCCD NET517 SKY130_FD_SC_HD__BUF_12
XINPUT518 MPRJ_ADR_O_CORE[10] VSSD VSSD VCCD VCCD NET518 SKY130_FD_SC_HD__CLKBUF_1
XINPUT519 MPRJ_ADR_O_CORE[11] VSSD VSSD VCCD VCCD NET519 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT52 LA_DATA_OUT_CORE[28] VSSD VSSD VCCD VCCD NET52 SKY130_FD_SC_HD__CLKBUF_4
XINPUT520 MPRJ_ADR_O_CORE[12] VSSD VSSD VCCD VCCD NET520 SKY130_FD_SC_HD__CLKBUF_2
XINPUT521 MPRJ_ADR_O_CORE[13] VSSD VSSD VCCD VCCD NET521 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT522 MPRJ_ADR_O_CORE[14] VSSD VSSD VCCD VCCD NET522 SKY130_FD_SC_HD__CLKBUF_2
XINPUT523 MPRJ_ADR_O_CORE[15] VSSD VSSD VCCD VCCD NET523 SKY130_FD_SC_HD__BUF_2
XINPUT524 MPRJ_ADR_O_CORE[16] VSSD VSSD VCCD VCCD NET524 SKY130_FD_SC_HD__BUF_2
XINPUT525 MPRJ_ADR_O_CORE[17] VSSD VSSD VCCD VCCD NET525 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT526 MPRJ_ADR_O_CORE[18] VSSD VSSD VCCD VCCD NET526 SKY130_FD_SC_HD__BUF_2
XINPUT527 MPRJ_ADR_O_CORE[19] VSSD VSSD VCCD VCCD NET527 SKY130_FD_SC_HD__CLKBUF_2
XINPUT528 MPRJ_ADR_O_CORE[1] VSSD VSSD VCCD VCCD NET528 SKY130_FD_SC_HD__CLKBUF_4
XINPUT529 MPRJ_ADR_O_CORE[20] VSSD VSSD VCCD VCCD NET529 SKY130_FD_SC_HD__CLKBUF_2
XINPUT53 LA_DATA_OUT_CORE[29] VSSD VSSD VCCD VCCD NET53 SKY130_FD_SC_HD__CLKBUF_4
XINPUT530 MPRJ_ADR_O_CORE[21] VSSD VSSD VCCD VCCD NET530 SKY130_FD_SC_HD__BUF_2
XINPUT531 MPRJ_ADR_O_CORE[22] VSSD VSSD VCCD VCCD NET531 SKY130_FD_SC_HD__CLKBUF_2
XINPUT532 MPRJ_ADR_O_CORE[23] VSSD VSSD VCCD VCCD NET532 SKY130_FD_SC_HD__CLKBUF_2
XINPUT533 MPRJ_ADR_O_CORE[24] VSSD VSSD VCCD VCCD NET533 SKY130_FD_SC_HD__CLKBUF_4
XINPUT534 MPRJ_ADR_O_CORE[25] VSSD VSSD VCCD VCCD NET534 SKY130_FD_SC_HD__BUF_2
XINPUT535 MPRJ_ADR_O_CORE[26] VSSD VSSD VCCD VCCD NET535 SKY130_FD_SC_HD__BUF_2
XINPUT536 MPRJ_ADR_O_CORE[27] VSSD VSSD VCCD VCCD NET536 SKY130_FD_SC_HD__BUF_2
XINPUT537 MPRJ_ADR_O_CORE[28] VSSD VSSD VCCD VCCD NET537 SKY130_FD_SC_HD__BUF_2
XINPUT538 MPRJ_ADR_O_CORE[29] VSSD VSSD VCCD VCCD NET538 SKY130_FD_SC_HD__BUF_2
XINPUT539 MPRJ_ADR_O_CORE[2] VSSD VSSD VCCD VCCD NET539 SKY130_FD_SC_HD__BUF_12
XINPUT54 LA_DATA_OUT_CORE[2] VSSD VSSD VCCD VCCD NET54 SKY130_FD_SC_HD__BUF_4
XINPUT540 MPRJ_ADR_O_CORE[30] VSSD VSSD VCCD VCCD NET540 SKY130_FD_SC_HD__BUF_2
XINPUT541 MPRJ_ADR_O_CORE[31] VSSD VSSD VCCD VCCD NET541 SKY130_FD_SC_HD__BUF_2
XINPUT542 MPRJ_ADR_O_CORE[3] VSSD VSSD VCCD VCCD NET542 SKY130_FD_SC_HD__CLKBUF_4
XINPUT543 MPRJ_ADR_O_CORE[4] VSSD VSSD VCCD VCCD NET543 SKY130_FD_SC_HD__BUF_12
XINPUT544 MPRJ_ADR_O_CORE[5] VSSD VSSD VCCD VCCD NET544 SKY130_FD_SC_HD__CLKBUF_4
XINPUT545 MPRJ_ADR_O_CORE[6] VSSD VSSD VCCD VCCD NET545 SKY130_FD_SC_HD__CLKBUF_2
XINPUT546 MPRJ_ADR_O_CORE[7] VSSD VSSD VCCD VCCD NET546 SKY130_FD_SC_HD__BUF_2
XINPUT547 MPRJ_ADR_O_CORE[8] VSSD VSSD VCCD VCCD NET547 SKY130_FD_SC_HD__BUF_2
XINPUT548 MPRJ_ADR_O_CORE[9] VSSD VSSD VCCD VCCD NET548 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT549 MPRJ_CYC_O_CORE VSSD VSSD VCCD VCCD NET549 SKY130_FD_SC_HD__CLKBUF_2
XINPUT55 LA_DATA_OUT_CORE[30] VSSD VSSD VCCD VCCD NET55 SKY130_FD_SC_HD__CLKBUF_4
XINPUT550 MPRJ_DAT_I_USER[0] VSSD VSSD VCCD VCCD NET550 SKY130_FD_SC_HD__BUF_12
XINPUT551 MPRJ_DAT_I_USER[10] VSSD VSSD VCCD VCCD NET551 SKY130_FD_SC_HD__BUF_12
XINPUT552 MPRJ_DAT_I_USER[11] VSSD VSSD VCCD VCCD NET552 SKY130_FD_SC_HD__BUF_12
XINPUT553 MPRJ_DAT_I_USER[12] VSSD VSSD VCCD VCCD NET553 SKY130_FD_SC_HD__BUF_12
XINPUT554 MPRJ_DAT_I_USER[13] VSSD VSSD VCCD VCCD NET554 SKY130_FD_SC_HD__BUF_12
XINPUT555 MPRJ_DAT_I_USER[14] VSSD VSSD VCCD VCCD NET555 SKY130_FD_SC_HD__BUF_12
XINPUT556 MPRJ_DAT_I_USER[15] VSSD VSSD VCCD VCCD NET556 SKY130_FD_SC_HD__BUF_12
XINPUT557 MPRJ_DAT_I_USER[16] VSSD VSSD VCCD VCCD NET557 SKY130_FD_SC_HD__BUF_12
XINPUT558 MPRJ_DAT_I_USER[17] VSSD VSSD VCCD VCCD NET558 SKY130_FD_SC_HD__BUF_12
XINPUT559 MPRJ_DAT_I_USER[18] VSSD VSSD VCCD VCCD NET559 SKY130_FD_SC_HD__BUF_12
XINPUT56 LA_DATA_OUT_CORE[31] VSSD VSSD VCCD VCCD NET56 SKY130_FD_SC_HD__CLKBUF_4
XINPUT560 MPRJ_DAT_I_USER[19] VSSD VSSD VCCD VCCD NET560 SKY130_FD_SC_HD__BUF_12
XINPUT561 MPRJ_DAT_I_USER[1] VSSD VSSD VCCD VCCD NET561 SKY130_FD_SC_HD__CLKBUF_16
XINPUT562 MPRJ_DAT_I_USER[20] VSSD VSSD VCCD VCCD NET562 SKY130_FD_SC_HD__CLKBUF_16
XINPUT563 MPRJ_DAT_I_USER[21] VSSD VSSD VCCD VCCD NET563 SKY130_FD_SC_HD__BUF_8
XINPUT564 MPRJ_DAT_I_USER[22] VSSD VSSD VCCD VCCD NET564 SKY130_FD_SC_HD__BUF_8
XINPUT565 MPRJ_DAT_I_USER[23] VSSD VSSD VCCD VCCD NET565 SKY130_FD_SC_HD__BUF_6
XINPUT566 MPRJ_DAT_I_USER[24] VSSD VSSD VCCD VCCD NET566 SKY130_FD_SC_HD__BUF_2
XINPUT567 MPRJ_DAT_I_USER[25] VSSD VSSD VCCD VCCD NET567 SKY130_FD_SC_HD__CLKBUF_2
XINPUT568 MPRJ_DAT_I_USER[26] VSSD VSSD VCCD VCCD NET568 SKY130_FD_SC_HD__CLKBUF_2
XINPUT569 MPRJ_DAT_I_USER[27] VSSD VSSD VCCD VCCD NET569 SKY130_FD_SC_HD__CLKBUF_2
XINPUT57 LA_DATA_OUT_CORE[32] VSSD VSSD VCCD VCCD NET57 SKY130_FD_SC_HD__BUF_4
XINPUT570 MPRJ_DAT_I_USER[28] VSSD VSSD VCCD VCCD NET570 SKY130_FD_SC_HD__CLKBUF_2
XINPUT571 MPRJ_DAT_I_USER[29] VSSD VSSD VCCD VCCD NET571 SKY130_FD_SC_HD__CLKBUF_2
XINPUT572 MPRJ_DAT_I_USER[2] VSSD VSSD VCCD VCCD NET572 SKY130_FD_SC_HD__BUF_8
XINPUT573 MPRJ_DAT_I_USER[30] VSSD VSSD VCCD VCCD NET573 SKY130_FD_SC_HD__CLKBUF_2
XINPUT574 MPRJ_DAT_I_USER[31] VSSD VSSD VCCD VCCD NET574 SKY130_FD_SC_HD__CLKBUF_2
XINPUT575 MPRJ_DAT_I_USER[3] VSSD VSSD VCCD VCCD NET575 SKY130_FD_SC_HD__BUF_8
XINPUT576 MPRJ_DAT_I_USER[4] VSSD VSSD VCCD VCCD NET576 SKY130_FD_SC_HD__CLKBUF_16
XINPUT577 MPRJ_DAT_I_USER[5] VSSD VSSD VCCD VCCD NET577 SKY130_FD_SC_HD__BUF_12
XINPUT578 MPRJ_DAT_I_USER[6] VSSD VSSD VCCD VCCD NET578 SKY130_FD_SC_HD__BUF_12
XINPUT579 MPRJ_DAT_I_USER[7] VSSD VSSD VCCD VCCD NET579 SKY130_FD_SC_HD__BUF_8
XINPUT58 LA_DATA_OUT_CORE[33] VSSD VSSD VCCD VCCD NET58 SKY130_FD_SC_HD__BUF_4
XINPUT580 MPRJ_DAT_I_USER[8] VSSD VSSD VCCD VCCD NET580 SKY130_FD_SC_HD__CLKBUF_16
XINPUT581 MPRJ_DAT_I_USER[9] VSSD VSSD VCCD VCCD NET581 SKY130_FD_SC_HD__CLKBUF_16
XINPUT582 MPRJ_DAT_O_CORE[0] VSSD VSSD VCCD VCCD NET582 SKY130_FD_SC_HD__CLKBUF_2
XINPUT583 MPRJ_DAT_O_CORE[10] VSSD VSSD VCCD VCCD NET583 SKY130_FD_SC_HD__CLKBUF_2
XINPUT584 MPRJ_DAT_O_CORE[11] VSSD VSSD VCCD VCCD NET584 SKY130_FD_SC_HD__BUF_2
XINPUT585 MPRJ_DAT_O_CORE[12] VSSD VSSD VCCD VCCD NET585 SKY130_FD_SC_HD__BUF_2
XINPUT586 MPRJ_DAT_O_CORE[13] VSSD VSSD VCCD VCCD NET586 SKY130_FD_SC_HD__CLKBUF_4
XINPUT587 MPRJ_DAT_O_CORE[14] VSSD VSSD VCCD VCCD NET587 SKY130_FD_SC_HD__CLKBUF_2
XINPUT588 MPRJ_DAT_O_CORE[15] VSSD VSSD VCCD VCCD NET588 SKY130_FD_SC_HD__CLKBUF_2
XINPUT589 MPRJ_DAT_O_CORE[16] VSSD VSSD VCCD VCCD NET589 SKY130_FD_SC_HD__CLKBUF_2
XINPUT59 LA_DATA_OUT_CORE[34] VSSD VSSD VCCD VCCD NET59 SKY130_FD_SC_HD__BUF_4
XINPUT590 MPRJ_DAT_O_CORE[17] VSSD VSSD VCCD VCCD NET590 SKY130_FD_SC_HD__CLKBUF_2
XINPUT591 MPRJ_DAT_O_CORE[18] VSSD VSSD VCCD VCCD NET591 SKY130_FD_SC_HD__CLKBUF_2
XINPUT592 MPRJ_DAT_O_CORE[19] VSSD VSSD VCCD VCCD NET592 SKY130_FD_SC_HD__CLKBUF_2
XINPUT593 MPRJ_DAT_O_CORE[1] VSSD VSSD VCCD VCCD NET593 SKY130_FD_SC_HD__CLKBUF_2
XINPUT594 MPRJ_DAT_O_CORE[20] VSSD VSSD VCCD VCCD NET594 SKY130_FD_SC_HD__CLKBUF_2
XINPUT595 MPRJ_DAT_O_CORE[21] VSSD VSSD VCCD VCCD NET595 SKY130_FD_SC_HD__BUF_2
XINPUT596 MPRJ_DAT_O_CORE[22] VSSD VSSD VCCD VCCD NET596 SKY130_FD_SC_HD__CLKBUF_2
XINPUT597 MPRJ_DAT_O_CORE[23] VSSD VSSD VCCD VCCD NET597 SKY130_FD_SC_HD__CLKBUF_2
XINPUT598 MPRJ_DAT_O_CORE[24] VSSD VSSD VCCD VCCD NET598 SKY130_FD_SC_HD__BUF_2
XINPUT599 MPRJ_DAT_O_CORE[25] VSSD VSSD VCCD VCCD NET599 SKY130_FD_SC_HD__CLKBUF_2
XINPUT6 LA_DATA_OUT_CORE[101] VSSD VSSD VCCD VCCD NET6 SKY130_FD_SC_HD__BUF_4
XINPUT60 LA_DATA_OUT_CORE[35] VSSD VSSD VCCD VCCD NET60 SKY130_FD_SC_HD__CLKBUF_4
XINPUT600 MPRJ_DAT_O_CORE[26] VSSD VSSD VCCD VCCD NET600 SKY130_FD_SC_HD__BUF_2
XINPUT601 MPRJ_DAT_O_CORE[27] VSSD VSSD VCCD VCCD NET601 SKY130_FD_SC_HD__CLKBUF_2
XINPUT602 MPRJ_DAT_O_CORE[28] VSSD VSSD VCCD VCCD NET602 SKY130_FD_SC_HD__CLKBUF_2
XINPUT603 MPRJ_DAT_O_CORE[29] VSSD VSSD VCCD VCCD NET603 SKY130_FD_SC_HD__CLKBUF_2
XINPUT604 MPRJ_DAT_O_CORE[2] VSSD VSSD VCCD VCCD NET604 SKY130_FD_SC_HD__CLKBUF_2
XINPUT605 MPRJ_DAT_O_CORE[30] VSSD VSSD VCCD VCCD NET605 SKY130_FD_SC_HD__CLKBUF_2
XINPUT606 MPRJ_DAT_O_CORE[31] VSSD VSSD VCCD VCCD NET606 SKY130_FD_SC_HD__CLKBUF_2
XINPUT607 MPRJ_DAT_O_CORE[3] VSSD VSSD VCCD VCCD NET607 SKY130_FD_SC_HD__CLKBUF_2
XINPUT608 MPRJ_DAT_O_CORE[4] VSSD VSSD VCCD VCCD NET608 SKY130_FD_SC_HD__CLKBUF_2
XINPUT609 MPRJ_DAT_O_CORE[5] VSSD VSSD VCCD VCCD NET609 SKY130_FD_SC_HD__CLKBUF_2
XINPUT61 LA_DATA_OUT_CORE[36] VSSD VSSD VCCD VCCD NET61 SKY130_FD_SC_HD__CLKBUF_4
XINPUT610 MPRJ_DAT_O_CORE[6] VSSD VSSD VCCD VCCD NET610 SKY130_FD_SC_HD__CLKBUF_2
XINPUT611 MPRJ_DAT_O_CORE[7] VSSD VSSD VCCD VCCD NET611 SKY130_FD_SC_HD__CLKBUF_2
XINPUT612 MPRJ_DAT_O_CORE[8] VSSD VSSD VCCD VCCD NET612 SKY130_FD_SC_HD__CLKBUF_2
XINPUT613 MPRJ_DAT_O_CORE[9] VSSD VSSD VCCD VCCD NET613 SKY130_FD_SC_HD__CLKBUF_2
XINPUT614 MPRJ_IENA_WB VSSD VSSD VCCD VCCD NET614 SKY130_FD_SC_HD__BUF_6
XINPUT615 MPRJ_SEL_O_CORE[0] VSSD VSSD VCCD VCCD NET615 SKY130_FD_SC_HD__DLYMETAL6S2S_1
XINPUT616 MPRJ_SEL_O_CORE[1] VSSD VSSD VCCD VCCD NET616 SKY130_FD_SC_HD__CLKBUF_2
XINPUT617 MPRJ_SEL_O_CORE[2] VSSD VSSD VCCD VCCD NET617 SKY130_FD_SC_HD__BUF_2
XINPUT618 MPRJ_SEL_O_CORE[3] VSSD VSSD VCCD VCCD NET618 SKY130_FD_SC_HD__CLKBUF_1
XINPUT619 MPRJ_STB_O_CORE VSSD VSSD VCCD VCCD NET619 SKY130_FD_SC_HD__CLKBUF_4
XINPUT62 LA_DATA_OUT_CORE[37] VSSD VSSD VCCD VCCD NET62 SKY130_FD_SC_HD__CLKBUF_4
XINPUT620 MPRJ_WE_O_CORE VSSD VSSD VCCD VCCD NET620 SKY130_FD_SC_HD__CLKBUF_2
XINPUT621 USER_IRQ_CORE[0] VSSD VSSD VCCD VCCD NET621 SKY130_FD_SC_HD__CLKBUF_1
XINPUT622 USER_IRQ_CORE[1] VSSD VSSD VCCD VCCD NET622 SKY130_FD_SC_HD__CLKBUF_1
XINPUT623 USER_IRQ_CORE[2] VSSD VSSD VCCD VCCD NET623 SKY130_FD_SC_HD__CLKBUF_1
XINPUT624 USER_IRQ_ENA[0] VSSD VSSD VCCD VCCD NET624 SKY130_FD_SC_HD__CLKBUF_1
XINPUT625 USER_IRQ_ENA[1] VSSD VSSD VCCD VCCD NET625 SKY130_FD_SC_HD__CLKBUF_1
XINPUT626 USER_IRQ_ENA[2] VSSD VSSD VCCD VCCD NET626 SKY130_FD_SC_HD__CLKBUF_1
XINPUT63 LA_DATA_OUT_CORE[38] VSSD VSSD VCCD VCCD NET63 SKY130_FD_SC_HD__CLKBUF_4
XINPUT64 LA_DATA_OUT_CORE[39] VSSD VSSD VCCD VCCD NET64 SKY130_FD_SC_HD__CLKBUF_4
XINPUT65 LA_DATA_OUT_CORE[3] VSSD VSSD VCCD VCCD NET65 SKY130_FD_SC_HD__BUF_4
XINPUT66 LA_DATA_OUT_CORE[40] VSSD VSSD VCCD VCCD NET66 SKY130_FD_SC_HD__CLKBUF_4
XINPUT67 LA_DATA_OUT_CORE[41] VSSD VSSD VCCD VCCD NET67 SKY130_FD_SC_HD__CLKBUF_4
XINPUT68 LA_DATA_OUT_CORE[42] VSSD VSSD VCCD VCCD NET68 SKY130_FD_SC_HD__CLKBUF_4
XINPUT69 LA_DATA_OUT_CORE[43] VSSD VSSD VCCD VCCD NET69 SKY130_FD_SC_HD__CLKBUF_4
XINPUT7 LA_DATA_OUT_CORE[102] VSSD VSSD VCCD VCCD NET7 SKY130_FD_SC_HD__BUF_4
XINPUT70 LA_DATA_OUT_CORE[44] VSSD VSSD VCCD VCCD NET70 SKY130_FD_SC_HD__CLKBUF_4
XINPUT71 LA_DATA_OUT_CORE[45] VSSD VSSD VCCD VCCD NET71 SKY130_FD_SC_HD__BUF_4
XINPUT72 LA_DATA_OUT_CORE[46] VSSD VSSD VCCD VCCD NET72 SKY130_FD_SC_HD__BUF_4
XINPUT73 LA_DATA_OUT_CORE[47] VSSD VSSD VCCD VCCD NET73 SKY130_FD_SC_HD__BUF_4
XINPUT74 LA_DATA_OUT_CORE[48] VSSD VSSD VCCD VCCD NET74 SKY130_FD_SC_HD__CLKBUF_4
XINPUT75 LA_DATA_OUT_CORE[49] VSSD VSSD VCCD VCCD NET75 SKY130_FD_SC_HD__BUF_4
XINPUT76 LA_DATA_OUT_CORE[4] VSSD VSSD VCCD VCCD NET76 SKY130_FD_SC_HD__BUF_4
XINPUT77 LA_DATA_OUT_CORE[50] VSSD VSSD VCCD VCCD NET77 SKY130_FD_SC_HD__BUF_4
XINPUT78 LA_DATA_OUT_CORE[51] VSSD VSSD VCCD VCCD NET78 SKY130_FD_SC_HD__BUF_4
XINPUT79 LA_DATA_OUT_CORE[52] VSSD VSSD VCCD VCCD NET79 SKY130_FD_SC_HD__BUF_4
XINPUT8 LA_DATA_OUT_CORE[103] VSSD VSSD VCCD VCCD NET8 SKY130_FD_SC_HD__BUF_4
XINPUT80 LA_DATA_OUT_CORE[53] VSSD VSSD VCCD VCCD NET80 SKY130_FD_SC_HD__BUF_4
XINPUT81 LA_DATA_OUT_CORE[54] VSSD VSSD VCCD VCCD NET81 SKY130_FD_SC_HD__CLKBUF_4
XINPUT82 LA_DATA_OUT_CORE[55] VSSD VSSD VCCD VCCD NET82 SKY130_FD_SC_HD__BUF_4
XINPUT83 LA_DATA_OUT_CORE[56] VSSD VSSD VCCD VCCD NET83 SKY130_FD_SC_HD__CLKBUF_4
XINPUT84 LA_DATA_OUT_CORE[57] VSSD VSSD VCCD VCCD NET84 SKY130_FD_SC_HD__BUF_4
XINPUT85 LA_DATA_OUT_CORE[58] VSSD VSSD VCCD VCCD NET85 SKY130_FD_SC_HD__BUF_4
XINPUT86 LA_DATA_OUT_CORE[59] VSSD VSSD VCCD VCCD NET86 SKY130_FD_SC_HD__BUF_4
XINPUT87 LA_DATA_OUT_CORE[5] VSSD VSSD VCCD VCCD NET87 SKY130_FD_SC_HD__BUF_4
XINPUT88 LA_DATA_OUT_CORE[60] VSSD VSSD VCCD VCCD NET88 SKY130_FD_SC_HD__BUF_4
XINPUT89 LA_DATA_OUT_CORE[61] VSSD VSSD VCCD VCCD NET89 SKY130_FD_SC_HD__BUF_4
XINPUT9 LA_DATA_OUT_CORE[104] VSSD VSSD VCCD VCCD NET9 SKY130_FD_SC_HD__CLKBUF_4
XINPUT90 LA_DATA_OUT_CORE[62] VSSD VSSD VCCD VCCD NET90 SKY130_FD_SC_HD__BUF_4
XINPUT91 LA_DATA_OUT_CORE[63] VSSD VSSD VCCD VCCD NET91 SKY130_FD_SC_HD__BUF_4
XINPUT92 LA_DATA_OUT_CORE[64] VSSD VSSD VCCD VCCD NET92 SKY130_FD_SC_HD__BUF_4
XINPUT93 LA_DATA_OUT_CORE[65] VSSD VSSD VCCD VCCD NET93 SKY130_FD_SC_HD__BUF_4
XINPUT94 LA_DATA_OUT_CORE[66] VSSD VSSD VCCD VCCD NET94 SKY130_FD_SC_HD__BUF_4
XINPUT95 LA_DATA_OUT_CORE[67] VSSD VSSD VCCD VCCD NET95 SKY130_FD_SC_HD__BUF_4
XINPUT96 LA_DATA_OUT_CORE[68] VSSD VSSD VCCD VCCD NET96 SKY130_FD_SC_HD__BUF_4
XINPUT97 LA_DATA_OUT_CORE[69] VSSD VSSD VCCD VCCD NET97 SKY130_FD_SC_HD__BUF_4
XINPUT98 LA_DATA_OUT_CORE[6] VSSD VSSD VCCD VCCD NET98 SKY130_FD_SC_HD__BUF_4
XINPUT99 LA_DATA_OUT_CORE[70] VSSD VSSD VCCD VCCD NET99 SKY130_FD_SC_HD__BUF_4
X\LA_BUF[0] _073_ \LA_DATA_OUT_ENABLE[0]  VSSD VSSD VCCD VCCD NET627 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[100] _074_ \LA_DATA_OUT_ENABLE[100]  VSSD VSSD VCCD VCCD NET628 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[101] _075_ \LA_DATA_OUT_ENABLE[101]  VSSD VSSD VCCD VCCD NET629 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[102] _076_ \LA_DATA_OUT_ENABLE[102]  VSSD VSSD VCCD VCCD NET630 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[103] _077_ \LA_DATA_OUT_ENABLE[103]  VSSD VSSD VCCD VCCD NET631 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[104] _078_ \LA_DATA_OUT_ENABLE[104]  VSSD VSSD VCCD VCCD NET632 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[105] _079_ \LA_DATA_OUT_ENABLE[105]  VSSD VSSD VCCD VCCD NET633 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[106] _080_ \LA_DATA_OUT_ENABLE[106]  VSSD VSSD VCCD VCCD NET634 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[107] _081_ \LA_DATA_OUT_ENABLE[107]  VSSD VSSD VCCD VCCD NET635 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[108] _082_ \LA_DATA_OUT_ENABLE[108]  VSSD VSSD VCCD VCCD NET636 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[109] _083_ \LA_DATA_OUT_ENABLE[109]  VSSD VSSD VCCD VCCD NET637 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[10] _084_ \LA_DATA_OUT_ENABLE[10]  VSSD VSSD VCCD VCCD NET638 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[110] _085_ \LA_DATA_OUT_ENABLE[110]  VSSD VSSD VCCD VCCD NET639 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[111] _086_ \LA_DATA_OUT_ENABLE[111]  VSSD VSSD VCCD VCCD NET640 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[112] _087_ \LA_DATA_OUT_ENABLE[112]  VSSD VSSD VCCD VCCD NET641 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[113] _088_ \LA_DATA_OUT_ENABLE[113]  VSSD VSSD VCCD VCCD NET642 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[114] _089_ \LA_DATA_OUT_ENABLE[114]  VSSD VSSD VCCD VCCD NET643 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[115] _090_ \LA_DATA_OUT_ENABLE[115]  VSSD VSSD VCCD VCCD NET644 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[116] _091_ \LA_DATA_OUT_ENABLE[116]  VSSD VSSD VCCD VCCD NET645 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[117] _092_ \LA_DATA_OUT_ENABLE[117]  VSSD VSSD VCCD VCCD NET646 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[118] _093_ \LA_DATA_OUT_ENABLE[118]  VSSD VSSD VCCD VCCD NET647 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[119] _094_ \LA_DATA_OUT_ENABLE[119]  VSSD VSSD VCCD VCCD NET648 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[11] _095_ \LA_DATA_OUT_ENABLE[11]  VSSD VSSD VCCD VCCD NET649 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[120] _096_ \LA_DATA_OUT_ENABLE[120]  VSSD VSSD VCCD VCCD NET650 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[121] _097_ \LA_DATA_OUT_ENABLE[121]  VSSD VSSD VCCD VCCD NET651 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[122] _098_ \LA_DATA_OUT_ENABLE[122]  VSSD VSSD VCCD VCCD NET652 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[123] _099_ \LA_DATA_OUT_ENABLE[123]  VSSD VSSD VCCD VCCD NET653 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[124] _100_ \LA_DATA_OUT_ENABLE[124]  VSSD VSSD VCCD VCCD NET654 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[125] _101_ \LA_DATA_OUT_ENABLE[125]  VSSD VSSD VCCD VCCD NET655 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[126] _102_ \LA_DATA_OUT_ENABLE[126]  VSSD VSSD VCCD VCCD NET656 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[127] _103_ \LA_DATA_OUT_ENABLE[127]  VSSD VSSD VCCD VCCD NET657 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[12] _104_ \LA_DATA_OUT_ENABLE[12]  VSSD VSSD VCCD VCCD NET658 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[13] _105_ \LA_DATA_OUT_ENABLE[13]  VSSD VSSD VCCD VCCD NET659 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[14] _106_ \LA_DATA_OUT_ENABLE[14]  VSSD VSSD VCCD VCCD NET660 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[15] _107_ \LA_DATA_OUT_ENABLE[15]  VSSD VSSD VCCD VCCD NET661 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[16] _108_ \LA_DATA_OUT_ENABLE[16]  VSSD VSSD VCCD VCCD NET662 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[17] _109_ \LA_DATA_OUT_ENABLE[17]  VSSD VSSD VCCD VCCD NET663 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[18] _110_ \LA_DATA_OUT_ENABLE[18]  VSSD VSSD VCCD VCCD NET664 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[19] _111_ \LA_DATA_OUT_ENABLE[19]  VSSD VSSD VCCD VCCD NET665 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[1] _112_ \LA_DATA_OUT_ENABLE[1]  VSSD VSSD VCCD VCCD NET666 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[20] _113_ \LA_DATA_OUT_ENABLE[20]  VSSD VSSD VCCD VCCD NET667 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[21] _114_ \LA_DATA_OUT_ENABLE[21]  VSSD VSSD VCCD VCCD NET668 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[22] _115_ \LA_DATA_OUT_ENABLE[22]  VSSD VSSD VCCD VCCD NET669 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[23] _116_ \LA_DATA_OUT_ENABLE[23]  VSSD VSSD VCCD VCCD NET670 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[24] _117_ \LA_DATA_OUT_ENABLE[24]  VSSD VSSD VCCD VCCD NET671 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[25] _118_ \LA_DATA_OUT_ENABLE[25]  VSSD VSSD VCCD VCCD NET672 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[26] _119_ \LA_DATA_OUT_ENABLE[26]  VSSD VSSD VCCD VCCD NET673 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[27] _120_ \LA_DATA_OUT_ENABLE[27]  VSSD VSSD VCCD VCCD NET674 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[28] _121_ \LA_DATA_OUT_ENABLE[28]  VSSD VSSD VCCD VCCD NET675 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[29] _122_ \LA_DATA_OUT_ENABLE[29]  VSSD VSSD VCCD VCCD NET676 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[2] _123_ \LA_DATA_OUT_ENABLE[2]  VSSD VSSD VCCD VCCD NET677 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[30] _124_ \LA_DATA_OUT_ENABLE[30]  VSSD VSSD VCCD VCCD NET678 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[31] _125_ \LA_DATA_OUT_ENABLE[31]  VSSD VSSD VCCD VCCD NET679 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[32] _126_ \LA_DATA_OUT_ENABLE[32]  VSSD VSSD VCCD VCCD NET680 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[33] _127_ \LA_DATA_OUT_ENABLE[33]  VSSD VSSD VCCD VCCD NET681 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[34] _128_ \LA_DATA_OUT_ENABLE[34]  VSSD VSSD VCCD VCCD NET682 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[35] _129_ \LA_DATA_OUT_ENABLE[35]  VSSD VSSD VCCD VCCD NET683 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[36] _130_ \LA_DATA_OUT_ENABLE[36]  VSSD VSSD VCCD VCCD NET684 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[37] _131_ \LA_DATA_OUT_ENABLE[37]  VSSD VSSD VCCD VCCD NET685 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[38] _132_ \LA_DATA_OUT_ENABLE[38]  VSSD VSSD VCCD VCCD NET686 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[39] _133_ \LA_DATA_OUT_ENABLE[39]  VSSD VSSD VCCD VCCD NET687 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[3] _134_ \LA_DATA_OUT_ENABLE[3]  VSSD VSSD VCCD VCCD NET688 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[40] _135_ \LA_DATA_OUT_ENABLE[40]  VSSD VSSD VCCD VCCD NET689 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[41] _136_ \LA_DATA_OUT_ENABLE[41]  VSSD VSSD VCCD VCCD NET690 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[42] _137_ \LA_DATA_OUT_ENABLE[42]  VSSD VSSD VCCD VCCD NET691 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[43] _138_ \LA_DATA_OUT_ENABLE[43]  VSSD VSSD VCCD VCCD NET692 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[44] _139_ \LA_DATA_OUT_ENABLE[44]  VSSD VSSD VCCD VCCD NET693 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[45] _140_ \LA_DATA_OUT_ENABLE[45]  VSSD VSSD VCCD VCCD NET694 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[46] _141_ \LA_DATA_OUT_ENABLE[46]  VSSD VSSD VCCD VCCD NET695 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[47] _142_ \LA_DATA_OUT_ENABLE[47]  VSSD VSSD VCCD VCCD NET696 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[48] _143_ \LA_DATA_OUT_ENABLE[48]  VSSD VSSD VCCD VCCD NET697 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[49] _144_ \LA_DATA_OUT_ENABLE[49]  VSSD VSSD VCCD VCCD NET698 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[4] _145_ \LA_DATA_OUT_ENABLE[4]  VSSD VSSD VCCD VCCD NET699 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[50] _146_ \LA_DATA_OUT_ENABLE[50]  VSSD VSSD VCCD VCCD NET700 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[51] _147_ \LA_DATA_OUT_ENABLE[51]  VSSD VSSD VCCD VCCD NET701 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[52] _148_ \LA_DATA_OUT_ENABLE[52]  VSSD VSSD VCCD VCCD NET702 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[53] _149_ \LA_DATA_OUT_ENABLE[53]  VSSD VSSD VCCD VCCD NET703 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[54] _150_ \LA_DATA_OUT_ENABLE[54]  VSSD VSSD VCCD VCCD NET704 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[55] _151_ \LA_DATA_OUT_ENABLE[55]  VSSD VSSD VCCD VCCD NET705 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[56] _152_ \LA_DATA_OUT_ENABLE[56]  VSSD VSSD VCCD VCCD NET706 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[57] _153_ \LA_DATA_OUT_ENABLE[57]  VSSD VSSD VCCD VCCD NET707 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[58] _154_ \LA_DATA_OUT_ENABLE[58]  VSSD VSSD VCCD VCCD NET708 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[59] _155_ \LA_DATA_OUT_ENABLE[59]  VSSD VSSD VCCD VCCD NET709 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[5] _156_ \LA_DATA_OUT_ENABLE[5]  VSSD VSSD VCCD VCCD NET710 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[60] _157_ \LA_DATA_OUT_ENABLE[60]  VSSD VSSD VCCD VCCD NET711 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[61] _158_ \LA_DATA_OUT_ENABLE[61]  VSSD VSSD VCCD VCCD NET712 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[62] _159_ \LA_DATA_OUT_ENABLE[62]  VSSD VSSD VCCD VCCD NET713 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[63] _160_ \LA_DATA_OUT_ENABLE[63]  VSSD VSSD VCCD VCCD NET714 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[64] _161_ \LA_DATA_OUT_ENABLE[64]  VSSD VSSD VCCD VCCD NET715 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[65] _162_ \LA_DATA_OUT_ENABLE[65]  VSSD VSSD VCCD VCCD NET716 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[66] _163_ \LA_DATA_OUT_ENABLE[66]  VSSD VSSD VCCD VCCD NET717 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[67] _164_ \LA_DATA_OUT_ENABLE[67]  VSSD VSSD VCCD VCCD NET718 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[68] _165_ \LA_DATA_OUT_ENABLE[68]  VSSD VSSD VCCD VCCD NET719 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[69] _166_ \LA_DATA_OUT_ENABLE[69]  VSSD VSSD VCCD VCCD NET720 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[6] _167_ \LA_DATA_OUT_ENABLE[6]  VSSD VSSD VCCD VCCD NET721 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[70] _168_ \LA_DATA_OUT_ENABLE[70]  VSSD VSSD VCCD VCCD NET722 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[71] _169_ \LA_DATA_OUT_ENABLE[71]  VSSD VSSD VCCD VCCD NET723 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[72] _170_ \LA_DATA_OUT_ENABLE[72]  VSSD VSSD VCCD VCCD NET724 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[73] _171_ \LA_DATA_OUT_ENABLE[73]  VSSD VSSD VCCD VCCD NET725 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[74] _172_ \LA_DATA_OUT_ENABLE[74]  VSSD VSSD VCCD VCCD NET726 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[75] _173_ \LA_DATA_OUT_ENABLE[75]  VSSD VSSD VCCD VCCD NET727 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[76] _174_ \LA_DATA_OUT_ENABLE[76]  VSSD VSSD VCCD VCCD NET728 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[77] _175_ \LA_DATA_OUT_ENABLE[77]  VSSD VSSD VCCD VCCD NET729 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[78] _176_ \LA_DATA_OUT_ENABLE[78]  VSSD VSSD VCCD VCCD NET730 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[79] _177_ \LA_DATA_OUT_ENABLE[79]  VSSD VSSD VCCD VCCD NET731 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[7] _178_ \LA_DATA_OUT_ENABLE[7]  VSSD VSSD VCCD VCCD NET732 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[80] _179_ \LA_DATA_OUT_ENABLE[80]  VSSD VSSD VCCD VCCD NET733 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[81] _180_ \LA_DATA_OUT_ENABLE[81]  VSSD VSSD VCCD VCCD NET734 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[82] _181_ \LA_DATA_OUT_ENABLE[82]  VSSD VSSD VCCD VCCD NET735 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[83] _182_ \LA_DATA_OUT_ENABLE[83]  VSSD VSSD VCCD VCCD NET736 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[84] _183_ \LA_DATA_OUT_ENABLE[84]  VSSD VSSD VCCD VCCD NET737 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[85] _184_ \LA_DATA_OUT_ENABLE[85]  VSSD VSSD VCCD VCCD NET738 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[86] _185_ \LA_DATA_OUT_ENABLE[86]  VSSD VSSD VCCD VCCD NET739 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[87] _186_ \LA_DATA_OUT_ENABLE[87]  VSSD VSSD VCCD VCCD NET740 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[88] _187_ \LA_DATA_OUT_ENABLE[88]  VSSD VSSD VCCD VCCD NET741 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[89] _188_ \LA_DATA_OUT_ENABLE[89]  VSSD VSSD VCCD VCCD NET742 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[8] _189_ \LA_DATA_OUT_ENABLE[8]  VSSD VSSD VCCD VCCD NET743 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[90] _190_ \LA_DATA_OUT_ENABLE[90]  VSSD VSSD VCCD VCCD NET744 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[91] _191_ \LA_DATA_OUT_ENABLE[91]  VSSD VSSD VCCD VCCD NET745 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[92] _192_ \LA_DATA_OUT_ENABLE[92]  VSSD VSSD VCCD VCCD NET746 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[93] _193_ \LA_DATA_OUT_ENABLE[93]  VSSD VSSD VCCD VCCD NET747 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[94] _194_ \LA_DATA_OUT_ENABLE[94]  VSSD VSSD VCCD VCCD NET748 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[95] _195_ \LA_DATA_OUT_ENABLE[95]  VSSD VSSD VCCD VCCD NET749 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[96] _196_ \LA_DATA_OUT_ENABLE[96]  VSSD VSSD VCCD VCCD NET750 SKY130_FD_SC_HD__EINVP_4
X\LA_BUF[97] _197_ \LA_DATA_OUT_ENABLE[97]  VSSD VSSD VCCD VCCD NET751 SKY130_FD_SC_HD__EINVP_2
X\LA_BUF[98] _198_ \LA_DATA_OUT_ENABLE[98]  VSSD VSSD VCCD VCCD NET752 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[99] _199_ \LA_DATA_OUT_ENABLE[99]  VSSD VSSD VCCD VCCD NET753 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF[9] _200_ \LA_DATA_OUT_ENABLE[9]  VSSD VSSD VCCD VCCD NET754 SKY130_FD_SC_HD__EINVP_8
X\LA_BUF_ENABLE[0] NET388 \MPRJ_LOGIC1[74]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[0]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[100] NET389 \MPRJ_LOGIC1[174]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[100]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[101] NET390 \MPRJ_LOGIC1[175]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[101]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[102] NET391 \MPRJ_LOGIC1[176]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[102]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[103] NET392 \MPRJ_LOGIC1[177]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[103]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[104] NET393 \MPRJ_LOGIC1[178]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[104]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[105] NET394 \MPRJ_LOGIC1[179]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[105]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[106] NET395 \MPRJ_LOGIC1[180]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[106]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[107] NET396 \MPRJ_LOGIC1[181]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[107]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[108] NET397 \MPRJ_LOGIC1[182]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[108]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[109] NET398 \MPRJ_LOGIC1[183]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[109]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[10] NET399 \MPRJ_LOGIC1[84]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[10]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[110] NET400 \MPRJ_LOGIC1[184]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[110]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[111] NET401 \MPRJ_LOGIC1[185]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[111]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[112] NET402 \MPRJ_LOGIC1[186]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[112]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[113] NET403 \MPRJ_LOGIC1[187]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[113]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[114] NET404 \MPRJ_LOGIC1[188]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[114]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[115] NET405 \MPRJ_LOGIC1[189]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[115]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[116] NET406 \MPRJ_LOGIC1[190]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[116]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[117] NET407 \MPRJ_LOGIC1[191]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[117]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[118] NET408 \MPRJ_LOGIC1[192]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[118]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[119] NET409 \MPRJ_LOGIC1[193]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[119]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[11] NET410 \MPRJ_LOGIC1[85]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[11]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[120] NET411 \MPRJ_LOGIC1[194]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[120]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[121] NET412 \MPRJ_LOGIC1[195]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[121]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[122] NET413 \MPRJ_LOGIC1[196]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[122]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[123] NET414 \MPRJ_LOGIC1[197]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[123]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[124] NET415 \MPRJ_LOGIC1[198]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[124]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[125] NET416 \MPRJ_LOGIC1[199]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[125]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[126] NET417 \MPRJ_LOGIC1[200]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[126]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[127] NET418 \MPRJ_LOGIC1[201]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[127]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[12] NET419 \MPRJ_LOGIC1[86]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[12]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[13] NET420 \MPRJ_LOGIC1[87]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[13]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[14] NET421 \MPRJ_LOGIC1[88]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[14]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[15] NET422 \MPRJ_LOGIC1[89]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[15]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[16] NET423 \MPRJ_LOGIC1[90]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[16]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[17] NET424 \MPRJ_LOGIC1[91]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[17]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[18] NET425 \MPRJ_LOGIC1[92]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[18]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[19] NET426 \MPRJ_LOGIC1[93]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[19]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[1] NET427 \MPRJ_LOGIC1[75]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[1]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[20] NET428 \MPRJ_LOGIC1[94]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[20]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[21] NET429 \MPRJ_LOGIC1[95]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[21]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[22] NET430 \MPRJ_LOGIC1[96]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[22]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[23] NET431 \MPRJ_LOGIC1[97]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[23]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[24] NET432 \MPRJ_LOGIC1[98]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[24]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[25] NET433 \MPRJ_LOGIC1[99]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[25]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[26] NET434 \MPRJ_LOGIC1[100]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[26]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[27] NET435 \MPRJ_LOGIC1[101]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[27]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[28] NET436 \MPRJ_LOGIC1[102]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[28]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[29] NET437 \MPRJ_LOGIC1[103]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[29]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[2] NET438 \MPRJ_LOGIC1[76]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[2]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[30] NET439 \MPRJ_LOGIC1[104]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[30]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[31] NET440 \MPRJ_LOGIC1[105]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[31]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[32] NET441 \MPRJ_LOGIC1[106]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[32]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[33] NET442 \MPRJ_LOGIC1[107]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[33]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[34] NET443 \MPRJ_LOGIC1[108]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[34]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[35] NET444 \MPRJ_LOGIC1[109]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[35]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[36] NET445 \MPRJ_LOGIC1[110]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[36]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[37] NET446 \MPRJ_LOGIC1[111]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[37]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[38] NET447 \MPRJ_LOGIC1[112]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[38]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[39] NET448 \MPRJ_LOGIC1[113]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[39]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[3] NET449 \MPRJ_LOGIC1[77]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[3]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[40] NET450 \MPRJ_LOGIC1[114]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[40]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[41] NET451 \MPRJ_LOGIC1[115]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[41]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[42] NET452 \MPRJ_LOGIC1[116]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[42]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[43] NET453 \MPRJ_LOGIC1[117]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[43]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[44] NET454 \MPRJ_LOGIC1[118]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[44]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[45] NET455 \MPRJ_LOGIC1[119]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[45]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[46] NET456 \MPRJ_LOGIC1[120]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[46]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[47] NET457 \MPRJ_LOGIC1[121]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[47]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[48] NET458 \MPRJ_LOGIC1[122]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[48]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[49] NET459 \MPRJ_LOGIC1[123]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[49]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[4] NET460 \MPRJ_LOGIC1[78]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[4]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[50] NET461 \MPRJ_LOGIC1[124]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[50]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[51] NET462 \MPRJ_LOGIC1[125]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[51]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[52] NET463 \MPRJ_LOGIC1[126]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[52]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[53] NET464 \MPRJ_LOGIC1[127]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[53]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[54] NET465 \MPRJ_LOGIC1[128]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[54]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[55] NET466 \MPRJ_LOGIC1[129]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[55]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[56] NET467 \MPRJ_LOGIC1[130]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[56]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[57] NET468 \MPRJ_LOGIC1[131]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[57]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[58] NET469 \MPRJ_LOGIC1[132]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[58]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[59] NET470 \MPRJ_LOGIC1[133]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[59]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[5] NET471 \MPRJ_LOGIC1[79]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[5]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[60] NET472 \MPRJ_LOGIC1[134]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[60]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[61] NET473 \MPRJ_LOGIC1[135]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[61]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[62] NET474 \MPRJ_LOGIC1[136]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[62]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[63] NET475 \MPRJ_LOGIC1[137]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[63]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[64] NET476 \MPRJ_LOGIC1[138]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[64]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[65] NET477 \MPRJ_LOGIC1[139]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[65]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[66] NET478 \MPRJ_LOGIC1[140]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[66]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[67] NET479 \MPRJ_LOGIC1[141]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[67]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[68] NET480 \MPRJ_LOGIC1[142]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[68]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[69] NET481 \MPRJ_LOGIC1[143]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[69]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[6] NET482 \MPRJ_LOGIC1[80]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[6]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[70] NET483 \MPRJ_LOGIC1[144]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[70]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[71] NET484 \MPRJ_LOGIC1[145]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[71]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[72] NET485 \MPRJ_LOGIC1[146]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[72]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[73] NET486 \MPRJ_LOGIC1[147]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[73]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[74] NET487 \MPRJ_LOGIC1[148]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[74]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[75] NET488 \MPRJ_LOGIC1[149]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[75]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[76] NET489 \MPRJ_LOGIC1[150]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[76]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[77] NET490 \MPRJ_LOGIC1[151]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[77]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[78] NET491 \MPRJ_LOGIC1[152]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[78]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[79] NET492 \MPRJ_LOGIC1[153]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[79]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[7] NET493 \MPRJ_LOGIC1[81]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[7]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[80] NET494 \MPRJ_LOGIC1[154]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[80]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[81] NET495 \MPRJ_LOGIC1[155]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[81]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[82] NET496 \MPRJ_LOGIC1[156]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[82]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[83] NET497 \MPRJ_LOGIC1[157]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[83]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[84] NET498 \MPRJ_LOGIC1[158]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[84]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[85] NET499 \MPRJ_LOGIC1[159]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[85]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[86] NET500 \MPRJ_LOGIC1[160]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[86]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[87] NET501 \MPRJ_LOGIC1[161]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[87]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[88] NET502 \MPRJ_LOGIC1[162]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[88]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[89] NET503 \MPRJ_LOGIC1[163]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[89]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[8] NET504 \MPRJ_LOGIC1[82]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[8]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[90] NET505 \MPRJ_LOGIC1[164]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[90]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[91] NET506 \MPRJ_LOGIC1[165]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[91]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[92] NET507 \MPRJ_LOGIC1[166]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[92]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[93] NET508 \MPRJ_LOGIC1[167]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[93]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[94] NET509 \MPRJ_LOGIC1[168]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[94]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[95] NET510 \MPRJ_LOGIC1[169]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[95]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[96] NET511 \MPRJ_LOGIC1[170]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[96]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[97] NET512 \MPRJ_LOGIC1[171]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[97]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[98] NET513 \MPRJ_LOGIC1[172]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[98]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[99] NET514 \MPRJ_LOGIC1[173]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[99]  SKY130_FD_SC_HD__AND2B_1
X\LA_BUF_ENABLE[9] NET515 \MPRJ_LOGIC1[83]  VSSD VSSD VCCD VCCD \LA_DATA_OUT_ENABLE[9]  SKY130_FD_SC_HD__AND2B_1
