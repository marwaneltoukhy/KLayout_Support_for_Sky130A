* Extracted by KLayout on : 19/01/2022 09:20

.SUBCKT caravel_clocking ext_clk_sel VPWR sel[0] sel[1] sel[2] pll_clk sel2[0]
+ pll_clk90 ext_clk sel2[1] resetb sel2[2] ext_reset core_clk user_clk
+ resetb_sync VGND
X$1 VGND \$21 \$15 \$2 \$102 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$2 VPWR \$2 VPWR \$33 VGND \$29 VGND sky130_fd_sc_hd__xnor2_1
X$3 VPWR \$23 VPWR VGND \$10 \$3 VGND sky130_fd_sc_hd__nand2_1
X$4 VPWR \$3 VPWR VGND \$11 \$4 \$57 VGND sky130_fd_sc_hd__nand3_1
X$5 VPWR VPWR VGND \$73 \$4 VGND sky130_fd_sc_hd__clkbuf_2
X$6 VPWR \$110 VPWR VGND \$4 \$93 \$92 VGND sky130_fd_sc_hd__nand3_1
X$7 VPWR \$101 VPWR VGND \$4 \$79 \$80 VGND sky130_fd_sc_hd__nand3_1
X$8 VPWR \$30 VPWR VGND \$40 \$4 \$57 VGND sky130_fd_sc_hd__nand3_1
X$9 VPWR \$131 VPWR VGND \$122 \$4 \$123 VGND sky130_fd_sc_hd__nand3_1
X$10 VPWR \$18 VGND VPWR \$5 VGND sky130_fd_sc_hd__clkbuf_1
X$11 VGND \$5 \$48 \$47 \$31 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$12 VPWR \$19 VPWR \$13 VGND \$6 VGND sky130_fd_sc_hd__xnor2_1
X$13 VPWR \$13 \$76 VGND \$81 VPWR \$6 VGND sky130_fd_sc_hd__nor3_1
X$14 VPWR \$13 VPWR \$118 VGND \$81 \$6 VGND sky130_fd_sc_hd__o21a_1
X$15 VPWR \$6 VGND VPWR \$106 VGND sky130_fd_sc_hd__dlygate4sd1_1
X$16 VPWR \$6 VGND VPWR \$38 VGND sky130_fd_sc_hd__clkbuf_1
X$17 VGND \$7 \$20 \$14 \$67 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$18 VPWR \$7 VPWR VGND \$73 \$29 \$80 VGND sky130_fd_sc_hd__nand3_1
X$19 VPWR \$8 \$33 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$20 VGND \$22 \$9 \$8 \$102 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$21 VPWR \$9 VGND VPWR \$53 VGND sky130_fd_sc_hd__dlygate4sd1_1
X$22 VPWR \$38 VGND VPWR \$9 VGND sky130_fd_sc_hd__dlygate4sd1_1
X$23 VPWR \$10 VPWR VGND \$58 \$63 VGND sky130_fd_sc_hd__nand2_1
X$24 VGND \$35 \$11 \$39 \$23 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$25 VPWR \$45 VGND \$40 VPWR \$11 VGND sky130_fd_sc_hd__nor2_1
X$26 VPWR \$16 \$11 VPWR \$24 VGND VGND sky130_fd_sc_hd__xor2_1
X$27 VGND \$69 \$11 \$40 \$12 VPWR VPWR VGND sky130_fd_sc_hd__nor3b_2
X$28 VPWR VGND VPWR \$42 \$12 VGND sky130_fd_sc_hd__inv_2
X$29 VPWR \$16 VGND \$12 VPWR \$40 VGND sky130_fd_sc_hd__nor2_1
X$30 VGND \$35 \$12 \$39 \$51 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$31 VPWR \$55 VPWR VGND \$45 \$12 VGND sky130_fd_sc_hd__nand2_1
X$32 VPWR \$25 VPWR \$12 VGND \$40 VGND sky130_fd_sc_hd__xnor2_1
X$33 VPWR VPWR VGND \$71 \$13 VGND sky130_fd_sc_hd__clkbuf_2
X$34 VGND \$14 \$15 \$21 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$35 VPWR \$98 VGND \$15 VPWR \$103 VGND sky130_fd_sc_hd__or2b_1
X$36 VPWR VGND \$15 VPWR \$71 VGND sky130_fd_sc_hd__clkbuf_4
X$37 VPWR \$15 VGND \$98 VPWR \$117 VGND sky130_fd_sc_hd__or2b_1
X$38 VGND \$98 \$39 \$15 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$39 VPWR \$15 VPWR \$116 VGND \$38 \$128 VGND sky130_fd_sc_hd__o21a_1
X$40 VPWR \$151 VGND \$15 VPWR \$128 VGND sky130_fd_sc_hd__nor2_1
X$41 VGND \$133 \$15 \$127 \$130 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$42 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$43 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$44 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$45 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$46 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$47 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$48 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$49 VPWR \$15 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$50 VPWR \$26 VPWR VGND \$58 \$17 VGND sky130_fd_sc_hd__nand2_1
X$51 VGND \$17 \$38 \$52 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$52 VGND \$35 \$47 \$60 \$18 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$53 VGND \$48 \$19 \$49 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$54 VGND \$35 \$29 \$60 \$20 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$55 VGND \$56 \$53 \$22 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$56 VGND \$59 \$81 \$24 \$69 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$57 VGND \$70 \$71 \$25 \$69 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$58 VPWR VPWR \$42 VGND \$58 \$51 \$26 VGND sky130_fd_sc_hd__o21ai_1
X$59 VGND \$43 ext_clk_sel VPWR VPWR VGND sky130_fd_sc_hd__dlymetal6s2s_1
X$60 VPWR ext_clk_sel VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$61 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$62 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$63 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$64 VPWR \$288 VPWR VGND \$256 \$271 VGND sky130_fd_sc_hd__nand2_1
X$65 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$66 VPWR resetb VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$67 VGND resetb \$35 VPWR VPWR VGND sky130_fd_sc_hd__buf_12
X$68 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$69 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$70 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$71 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$72 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$73 VGND \$263 \$215 \$285 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$74 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$75 VPWR \$289 VPWR VGND \$252 \$286 \$197 VGND sky130_fd_sc_hd__nand3_1
X$76 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$77 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$79 VPWR VPWR VGND \$242 \$189 VGND sky130_fd_sc_hd__clkbuf_2
X$80 VPWR \$278 VPWR VGND \$246 \$221 \$216 VGND sky130_fd_sc_hd__nand3_1
X$81 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$82 VGND \$278 \$253 \$244 \$227 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$83 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$84 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$85 VGND \$279 \$290 \$287 \$227 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$86 VPWR \$279 VPWR VGND \$264 \$281 \$216 VGND sky130_fd_sc_hd__nand3_1
X$87 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$88 VGND \$287 \$215 \$282 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$89 VPWR \$260 VGND \$213 VPWR \$246 VGND sky130_fd_sc_hd__nor2_1
X$90 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$91 VGND \$282 \$215 \$261 \$230 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$92 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$93 VGND \$291 \$188 \$259 \$292 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$94 VPWR \$280 VPWR VGND \$283 \$281 \$277 VGND sky130_fd_sc_hd__nand3_1
X$95 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$96 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$97 VGND \$35 \$267 \$168 \$280 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$98 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$99 VPWR \$294 VGND \$190 VPWR \$215 VGND sky130_fd_sc_hd__nor2_1
X$100 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$101 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$102 VGND \$35 \$215 \$188 \$293 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$103 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$104 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$105 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$106 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$107 VGND \$35 \$304 \$297 \$298 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$108 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$109 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$110 VPWR \$307 VPWR VGND \$299 \$281 \$220 VGND sky130_fd_sc_hd__nand3_1
X$111 VGND \$252 \$299 \$304 \$233 VPWR VPWR VGND sky130_fd_sc_hd__nor3b_2
X$112 VPWR \$305 VGND \$304 VPWR \$299 VGND sky130_fd_sc_hd__nor2_1
X$113 VPWR \$295 VPWR VGND \$305 \$233 VGND sky130_fd_sc_hd__nand2_1
X$114 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$116 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$117 VGND \$285 \$215 \$321 \$252 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$118 VPWR VPWR \$295 VGND \$220 \$306 \$286 VGND sky130_fd_sc_hd__o21bai_1
X$119 VPWR \$308 VPWR VGND \$281 \$306 \$289 VGND sky130_fd_sc_hd__nand3_1
X$120 VPWR VGND VPWR \$286 \$300 VGND sky130_fd_sc_hd__inv_2
X$121 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$122 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$123 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$124 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$125 VGND \$35 \$264 \$189 \$290 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$126 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$127 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$128 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$129 VPWR ext_clk VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$130 VGND ext_clk \$309 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$131 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$132 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$133 VPWR VPWR VGND \$309 \$276 VGND sky130_fd_sc_hd__clkbuf_2
X$134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$135 VGND \$35 \$293 \$188 \$296 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$136 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$138 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$139 VGND \$35 \$303 \$301 \$302 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$140 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$141 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$142 VPWR \$303 \$310 VGND VPWR VGND sky130_fd_sc_hd__clkdlybuf4s25_1
X$143 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$145 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$147 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$148 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$149 VPWR \$104 VGND VPWR \$95 VGND sky130_fd_sc_hd__clkbuf_1
X$150 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$151 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$152 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$153 VPWR \$99 \$96 VPWR \$105 VGND VGND sky130_fd_sc_hd__xor2_1
X$154 VPWR \$88 VPWR \$47 VGND \$44 VGND sky130_fd_sc_hd__xnor2_1
X$155 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$156 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$157 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$158 VGND \$64 \$81 \$71 \$38 \$85 VPWR VPWR VGND sky130_fd_sc_hd__o211a_1
X$159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$160 VPWR \$71 VGND VPWR \$78 VGND sky130_fd_sc_hd__dlygate4sd1_1
X$161 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$162 VGND \$101 \$107 \$100 \$67 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$163 VGND \$108 \$54 \$72 \$102 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$164 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$165 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$167 VPWR VGND \$89 \$102 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$168 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$169 VPWR \$109 VGND VPWR \$38 VGND sky130_fd_sc_hd__clkbuf_1
X$170 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$171 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$172 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$173 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$174 VPWR \$92 VPWR VGND \$69 \$82 \$97 VGND sky130_fd_sc_hd__nand3_1
X$175 VPWR VGND VPWR \$82 \$112 VGND sky130_fd_sc_hd__inv_2
X$176 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$177 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$178 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$179 VGND \$35 \$32 \$39 \$94 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$180 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$181 VPWR \$111 VGND VPWR sel[0] VGND sky130_fd_sc_hd__clkbuf_1
X$182 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$183 VPWR \$74 VPWR VGND \$90 \$117 \$103 VGND sky130_fd_sc_hd__nand3_1
X$184 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$185 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$186 VGND \$35 \$96 \$60 \$104 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$187 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$188 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$189 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$190 VGND \$95 \$113 \$96 \$31 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$191 VGND \$113 \$118 \$105 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$192 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$193 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$194 VPWR \$77 VGND VPWR \$54 VGND sky130_fd_sc_hd__clkbuf_1
X$195 VGND \$35 \$79 \$60 \$107 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$196 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$197 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$198 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$199 VPWR VPWR \$80 VGND \$89 \$122 \$114 VGND sky130_fd_sc_hd__o21bai_1
X$200 VPWR \$123 \$89 VGND \$116 \$114 VPWR VGND sky130_fd_sc_hd__nand3b_1
X$201 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$202 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$203 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$204 VPWR VGND VPWR \$114 \$119 VGND sky130_fd_sc_hd__inv_2
X$205 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$206 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$207 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$208 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$209 VGND \$35 \$112 \$120 \$110 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$210 VPWR VPWR \$124 VGND \$115 \$83 \$116 VGND sky130_fd_sc_hd__o21ai_1
X$211 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$212 VPWR \$128 \$115 VPWR \$121 VGND VGND sky130_fd_sc_hd__and2_1
X$213 VGND \$35 \$125 \$138 \$111 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$214 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$215 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$216 VPWR sel[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$217 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$218 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$219 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$220 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$221 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$222 VPWR VGND VPWR \$60 \$36 VGND sky130_fd_sc_hd__inv_4
X$223 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$224 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$225 VPWR \$49 \$47 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$226 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$227 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$228 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$229 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$230 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$231 VGND \$31 \$67 \$32 \$64 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$232 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$233 VPWR \$65 VGND \$33 VPWR \$29 VGND sky130_fd_sc_hd__nor2_1
X$234 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$235 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$236 VGND \$66 \$61 \$56 \$67 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$237 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$238 VPWR VPWR VGND \$62 \$80 VGND sky130_fd_sc_hd__clkbuf_2
X$239 VPWR \$58 VPWR VGND \$57 \$73 VGND sky130_fd_sc_hd__nand2_1
X$240 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$241 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$242 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$243 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$244 VGND \$63 \$54 \$59 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$246 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$247 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$248 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$249 VPWR \$46 VPWR VGND \$58 \$68 VGND sky130_fd_sc_hd__nand2_1
X$250 VPWR VGND VPWR \$39 \$41 VGND sky130_fd_sc_hd__inv_4
X$251 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$252 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$253 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$254 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$255 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$256 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$257 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$258 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$259 VPWR \$37 VGND VPWR \$75 VGND sky130_fd_sc_hd__clkbuf_1
X$260 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$261 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$262 VPWR \$99 VGND \$47 VPWR \$44 VGND sky130_fd_sc_hd__nor2_1
X$263 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$264 VGND \$75 \$87 \$44 \$31 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$265 VGND \$87 \$84 \$88 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$266 VPWR \$84 VGND \$118 VPWR \$76 VGND sky130_fd_sc_hd__nor2_1
X$267 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$268 VGND \$77 \$78 \$85 \$50 VPWR \$57 VPWR VGND sky130_fd_sc_hd__o211ai_4
X$269 VPWR \$65 \$79 VPWR \$72 VGND VGND sky130_fd_sc_hd__xor2_1
X$270 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$271 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$272 VPWR \$66 VPWR VGND \$73 \$33 \$80 VGND sky130_fd_sc_hd__nand3_1
X$273 VPWR \$86 VGND \$29 VPWR \$79 VGND sky130_fd_sc_hd__nor2_1
X$274 VPWR \$89 VPWR VGND \$86 \$33 VGND sky130_fd_sc_hd__nand2_1
X$275 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$276 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$277 VPWR VPWR \$81 VGND \$71 \$62 \$38 VGND sky130_fd_sc_hd__o21ai_1
X$278 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$279 VPWR VGND \$32 \$73 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$280 VPWR VPWR \$67 \$73 VGND \$62 VGND sky130_fd_sc_hd__nand2_2
X$281 VPWR VPWR \$55 VGND \$57 \$93 \$82 VGND sky130_fd_sc_hd__o21bai_1
X$282 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$283 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$284 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$285 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$286 VPWR \$83 VPWR \$94 VGND \$67 \$74 VGND sky130_fd_sc_hd__o21a_1
X$287 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$288 VGND \$68 \$71 \$70 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$289 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$290 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$291 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$292 VGND \$90 \$39 \$38 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$293 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$294 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$295 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$296 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$297 VGND \$35 \$202 \$189 \$201 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$298 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$299 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$300 VPWR VGND VPWR \$189 \$183 VGND sky130_fd_sc_hd__inv_4
X$301 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$302 VGND \$35 \$164 \$183 \$174 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$303 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$304 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$305 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$306 VPWR \$203 VGND \$158 VPWR \$164 VGND sky130_fd_sc_hd__nor2_1
X$307 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$308 VGND \$176 \$204 \$175 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$309 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$310 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$311 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$312 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$313 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$314 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$315 VPWR \$190 VPWR \$205 VGND \$215 \$196 VGND sky130_fd_sc_hd__o21a_1
X$316 VGND \$35 \$158 \$189 \$177 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$317 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$318 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$319 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$320 VGND \$170 \$195 \$227 \$197 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$321 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$322 VPWR \$193 VPWR \$190 VGND \$196 VGND sky130_fd_sc_hd__xnor2_1
X$323 VGND \$178 \$193 \$171 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$324 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$325 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$326 VGND \$194 \$189 \$190 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$327 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$328 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$329 VPWR \$199 VPWR \$206 VGND \$227 \$157 VGND sky130_fd_sc_hd__o21a_1
X$330 VPWR \$190 VGND \$194 VPWR \$159 VGND sky130_fd_sc_hd__or2b_1
X$331 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$332 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$333 VPWR \$194 VGND \$190 VPWR \$166 VGND sky130_fd_sc_hd__or2b_1
X$334 VGND pll_clk \$172 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$335 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$336 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$337 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$338 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$339 VPWR pll_clk VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$340 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$341 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$342 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$344 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$345 VGND \$35 \$180 \$168 \$185 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$346 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$347 VPWR \$185 VGND VPWR \$200 VGND sky130_fd_sc_hd__clkbuf_1
X$348 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$350 VGND \$200 \$180 \$207 \$196 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$351 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$352 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$353 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$354 VPWR \$181 VPWR \$186 VGND \$180 VGND sky130_fd_sc_hd__xnor2_1
X$355 VGND \$207 \$215 \$181 \$198 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$356 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$357 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$358 VGND \$182 \$186 \$187 \$196 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$359 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$360 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$361 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$362 VPWR \$208 \$186 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$363 VGND \$35 \$169 \$168 \$162 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$364 VPWR \$161 VGND VPWR \$182 VGND sky130_fd_sc_hd__clkbuf_1
X$365 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$366 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$367 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$368 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$369 VPWR \$186 \$163 VGND \$196 VPWR \$180 VGND sky130_fd_sc_hd__nor3_1
X$370 VGND \$35 \$191 \$188 \$192 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$371 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$372 VGND \$198 \$180 \$169 \$186 VPWR VPWR VGND sky130_fd_sc_hd__nor3b_2
X$373 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$374 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$375 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$376 VPWR sel[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$377 VPWR \$139 VGND VPWR sel[2] VGND sky130_fd_sc_hd__clkbuf_1
X$378 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$379 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$380 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$381 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$382 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$383 VGND \$35 \$233 \$189 \$255 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$384 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$385 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$386 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$387 VPWR VPWR \$241 VGND \$256 \$255 \$243 VGND sky130_fd_sc_hd__o21ai_1
X$388 VGND \$234 \$196 \$245 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$389 VPWR \$270 VPWR VGND \$256 \$263 VGND sky130_fd_sc_hd__nand2_1
X$390 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$391 VPWR \$258 VPWR \$233 VGND \$304 VGND sky130_fd_sc_hd__xnor2_1
X$392 VGND \$245 \$196 \$241 \$252 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$393 VGND \$271 \$190 \$272 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$394 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$395 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$396 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$397 VGND \$272 \$190 \$258 \$252 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$398 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$399 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$400 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$401 VPWR \$256 VPWR VGND \$220 \$221 VGND sky130_fd_sc_hd__nand2_1
X$402 VPWR VGND \$195 \$221 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$403 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$404 VPWR VPWR \$215 VGND \$190 \$235 \$196 VGND sky130_fd_sc_hd__o21ai_1
X$405 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$406 VPWR VPWR VGND \$221 \$281 VGND sky130_fd_sc_hd__clkbuf_2
X$407 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$408 VGND \$35 \$246 \$189 \$253 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$409 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$410 VPWR \$260 \$264 VPWR \$261 VGND VGND sky130_fd_sc_hd__xor2_1
X$411 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$412 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$413 VGND \$273 \$60 \$269 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$414 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$415 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$416 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$417 VGND pll_clk90 \$242 VPWR VPWR VGND sky130_fd_sc_hd__clkbuf_16
X$418 VPWR \$248 VPWR \$213 VGND \$246 VGND sky130_fd_sc_hd__xnor2_1
X$419 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$420 VPWR \$273 \$274 VGND VPWR VGND sky130_fd_sc_hd__clkdlybuf4s25_1
X$421 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$422 VGND \$259 \$275 \$276 \$179 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$423 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$424 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$425 VGND \$236 \$190 \$248 \$230 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$426 VPWR VGND \$265 \$230 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$427 VPWR \$265 VPWR VGND \$249 \$213 VGND sky130_fd_sc_hd__nand2_1
X$428 VPWR pll_clk90 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$429 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$430 VPWR \$249 VGND \$246 VPWR \$264 VGND sky130_fd_sc_hd__nor2_1
X$431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$432 VPWR \$277 \$265 VGND \$231 \$266 VPWR VGND sky130_fd_sc_hd__nand3b_1
X$433 VPWR \$190 VPWR \$231 VGND \$196 \$215 VGND sky130_fd_sc_hd__o21a_1
X$434 VPWR VPWR \$216 VGND \$265 \$283 \$266 VGND sky130_fd_sc_hd__o21bai_1
X$435 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$436 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$437 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$438 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$439 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$440 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$441 VPWR \$250 VPWR \$300 VGND \$267 VGND sky130_fd_sc_hd__xnor2_1
X$442 VPWR VGND \$196 \$218 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$443 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$444 VGND \$218 \$251 \$188 \$216 \$250 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2ai_2
X$445 VPWR VGND VPWR \$266 \$267 VGND sky130_fd_sc_hd__inv_2
X$446 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$447 VGND \$35 \$254 \$188 \$262 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$448 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$450 VGND \$35 \$190 \$188 \$254 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_4
X$451 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$452 VGND \$251 \$168 \$240 \$294 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$453 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$454 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$455 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$456 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$457 VPWR sel2[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$458 VPWR \$262 VGND VPWR sel2[1] VGND sky130_fd_sc_hd__clkbuf_1
X$459 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$460 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$461 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$462 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$463 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$464 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$465 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$466 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$467 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$468 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$469 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$470 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$471 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$472 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$473 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$474 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$475 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$476 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$477 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$478 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$479 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$480 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$481 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$482 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$483 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$484 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$485 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$486 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$487 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$488 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$489 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$490 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$491 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$492 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$493 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$494 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$495 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$496 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$497 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$498 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$499 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$500 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$501 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$502 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$503 VGND \$35 \$44 \$36 \$37 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$504 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$505 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$506 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$507 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$508 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$509 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$510 VPWR \$50 VGND VPWR \$38 VGND sky130_fd_sc_hd__clkbuf_1
X$511 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$512 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$513 VGND \$35 \$33 \$39 \$61 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$514 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$515 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$516 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$517 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$518 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$519 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$520 VPWR \$34 VPWR VGND \$46 \$30 VGND sky130_fd_sc_hd__nand2_1
X$521 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$522 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$523 VGND \$35 \$40 \$41 \$34 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$524 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$525 VGND \$52 \$38 \$42 \$69 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$527 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$528 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$529 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$530 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$531 VPWR \$148 VGND VPWR \$136 VGND sky130_fd_sc_hd__clkbuf_1
X$532 VPWR \$174 VGND VPWR \$155 VGND sky130_fd_sc_hd__clkbuf_1
X$533 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$534 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$536 VGND \$35 \$142 \$60 \$148 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$537 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$538 VPWR \$175 VPWR \$158 VGND \$164 VGND sky130_fd_sc_hd__xnor2_1
X$539 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$540 VGND \$155 \$176 \$164 \$170 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$541 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$542 VPWR \$156 VPWR \$140 VGND \$142 VGND sky130_fd_sc_hd__xnor2_1
X$543 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$544 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$545 VGND \$144 \$128 \$156 \$130 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$546 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$547 VPWR \$130 VGND \$142 \$143 VPWR \$140 VGND sky130_fd_sc_hd__nor3b_1
X$548 VPWR \$177 VGND VPWR \$165 VGND sky130_fd_sc_hd__clkbuf_1
X$549 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$550 VGND \$165 \$178 \$158 \$170 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$551 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$552 VPWR \$145 \$143 VPWR \$149 VGND VGND sky130_fd_sc_hd__xor2_1
X$553 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$554 VPWR \$171 \$158 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$555 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$556 VGND \$35 \$143 \$60 \$149 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$557 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$558 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$559 VPWR VPWR VGND \$172 \$60 VGND sky130_fd_sc_hd__clkbuf_2
X$560 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$561 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$562 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$563 VPWR \$153 VPWR VGND \$140 \$137 \$146 VGND sky130_fd_sc_hd__nand3_1
X$564 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$565 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$566 VPWR \$150 VPWR \$153 VGND \$154 VGND sky130_fd_sc_hd__xnor2_1
X$567 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$568 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$569 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$570 VGND \$35 \$154 \$39 \$150 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$571 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$572 VPWR \$157 VPWR VGND \$167 \$159 \$166 VGND sky130_fd_sc_hd__nand3_1
X$573 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$574 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$575 VGND \$167 \$168 \$196 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$576 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$577 VGND \$141 \$39 \$154 \$151 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$578 VPWR VPWR VGND \$172 \$39 VGND sky130_fd_sc_hd__clkbuf_2
X$579 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$580 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$581 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$582 VGND \$35 \$179 \$39 \$160 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$583 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$584 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$585 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$586 VGND \$35 \$81 \$138 \$147 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$588 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$589 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$590 VGND \$35 \$186 \$168 \$161 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$591 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$592 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$593 VGND \$35 \$71 \$138 \$152 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_4
X$594 VPWR VPWR VGND \$81 \$54 VGND sky130_fd_sc_hd__clkbuf_2
X$595 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$596 VPWR \$163 \$169 VPWR \$162 VGND VGND sky130_fd_sc_hd__xor2_1
X$597 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$598 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$599 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$600 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$601 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$602 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$603 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$604 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$605 VPWR VGND VPWR \$189 \$297 VGND sky130_fd_sc_hd__inv_4
X$606 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$607 VPWR \$298 VPWR VGND \$288 \$311 VGND sky130_fd_sc_hd__nand2_1
X$608 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$609 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$610 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$611 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$612 VPWR \$311 VPWR VGND \$304 \$281 \$220 VGND sky130_fd_sc_hd__nand3_1
X$613 VGND \$35 \$299 \$189 \$313 VPWR VPWR VGND sky130_fd_sc_hd__dfrtn_1
X$614 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$615 VPWR \$313 VPWR VGND \$270 \$307 VGND sky130_fd_sc_hd__nand2_1
X$616 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$617 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$618 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$619 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$620 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$621 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$622 VPWR \$318 VGND \$233 VPWR \$304 VGND sky130_fd_sc_hd__nor2_1
X$623 VPWR \$318 \$299 VPWR \$321 VGND VGND sky130_fd_sc_hd__xor2_1
X$624 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$625 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$627 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$628 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$629 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$630 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$631 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$632 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$633 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$634 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$635 VGND \$35 \$300 \$314 \$308 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$636 VPWR VGND VPWR \$189 \$314 VGND sky130_fd_sc_hd__inv_4
X$637 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$638 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$639 VPWR core_clk VGND VPWR \$322 VGND sky130_fd_sc_hd__clkbuf_1
X$640 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$641 VPWR \$269 VGND VPWR \$323 VGND sky130_fd_sc_hd__buf_1
X$642 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$643 VPWR VPWR VGND \$309 \$328 VGND sky130_fd_sc_hd__clkbuf_2
X$644 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$645 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$646 VGND \$323 \$273 \$328 \$35 VPWR VPWR VGND sky130_fd_sc_hd__mux2_2
X$647 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$648 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$649 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$650 VGND \$35 \$275 \$39 \$274 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$651 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$652 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$653 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$654 VPWR user_clk VGND VPWR \$291 VGND sky130_fd_sc_hd__clkbuf_1
X$655 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$656 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$657 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$658 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$659 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$660 VGND \$35 \$292 \$39 \$179 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$661 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$662 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$663 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$664 VGND \$322 \$138 \$259 \$292 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$665 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$666 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$667 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$668 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$669 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$670 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$671 VGND \$35 \$319 \$315 \$316 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$672 VPWR VGND VPWR \$322 \$315 VGND sky130_fd_sc_hd__inv_4
X$673 VPWR VGND resetb_sync VPWR \$324 VGND sky130_fd_sc_hd__buf_2
X$674 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$675 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$676 VPWR VPWR VGND \$316 VGND sky130_fd_sc_hd__conb_1
X$677 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$678 VPWR VGND VPWR \$322 \$301 VGND sky130_fd_sc_hd__inv_4
X$679 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$680 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$681 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$682 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$683 VPWR \$319 \$302 VGND VPWR VGND sky130_fd_sc_hd__clkdlybuf4s25_1
X$684 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$685 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$686 VGND \$35 \$320 \$317 \$310 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$687 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$688 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$689 VPWR VGND VPWR \$322 \$317 VGND sky130_fd_sc_hd__inv_4
X$690 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$691 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$692 VPWR ext_reset VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$693 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$694 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$695 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$696 VPWR \$324 VGND \$320 VPWR \$326 VGND sky130_fd_sc_hd__nor2_1
X$697 VPWR sel2[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$698 VPWR \$326 VGND VPWR ext_reset VGND sky130_fd_sc_hd__clkbuf_1
X$699 VPWR \$296 VGND VPWR sel2[2] VGND sky130_fd_sc_hd__clkbuf_1
X$700 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$701 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$702 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$703 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$704 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$705 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$706 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$707 VPWR \$201 VGND VPWR \$209 VGND sky130_fd_sc_hd__clkbuf_1
X$708 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$709 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$710 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$711 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$712 VGND \$209 \$210 \$202 \$170 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$713 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$714 VPWR VGND VPWR \$241 \$233 VGND sky130_fd_sc_hd__inv_2
X$715 VPWR \$243 VPWR VGND \$256 \$234 VGND sky130_fd_sc_hd__nand2_1
X$716 VPWR \$211 VGND \$164 VPWR \$202 VGND sky130_fd_sc_hd__nor2_1
X$717 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$718 VPWR \$203 \$202 VPWR \$212 VGND VGND sky130_fd_sc_hd__xor2_1
X$719 VGND \$210 \$205 \$212 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$720 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$721 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$722 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$723 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$724 VGND \$215 \$190 \$211 \$196 VPWR \$220 VPWR VGND
+ sky130_fd_sc_hd__o211ai_4
X$725 VPWR \$190 \$226 VGND \$215 VPWR \$196 VGND sky130_fd_sc_hd__nor3_1
X$726 VPWR \$204 VGND \$205 VPWR \$226 VGND sky130_fd_sc_hd__nor2_1
X$727 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$728 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$729 VGND \$197 \$215 \$190 \$196 \$211 VPWR VPWR VGND sky130_fd_sc_hd__o211a_1
X$730 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$731 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$732 VPWR VPWR \$227 \$221 VGND \$235 VGND sky130_fd_sc_hd__nand2_2
X$733 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$734 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$735 VPWR \$222 VPWR VGND \$213 \$221 \$216 VGND sky130_fd_sc_hd__nand3_1
X$736 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$737 VGND \$35 \$213 \$168 \$223 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$738 VGND \$222 \$223 \$229 \$227 VPWR VPWR VGND sky130_fd_sc_hd__a21bo_1
X$739 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$740 VPWR VPWR VGND \$235 \$216 VGND sky130_fd_sc_hd__clkbuf_2
X$741 VGND \$229 \$196 \$228 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$742 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$743 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$744 VGND \$244 \$190 \$236 \$195 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$745 VGND \$35 \$195 \$168 \$206 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$746 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$747 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$748 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$749 VGND \$228 \$196 \$237 \$230 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$750 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$751 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$752 VGND \$214 \$168 \$215 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$753 VPWR \$237 \$213 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$754 VPWR VPWR VGND \$242 \$168 VGND sky130_fd_sc_hd__clkbuf_2
X$755 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$756 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$757 VPWR VPWR \$238 VGND \$224 \$199 \$231 VGND sky130_fd_sc_hd__o21ai_1
X$758 VPWR \$215 \$224 VPWR \$214 VGND VGND sky130_fd_sc_hd__and2_1
X$759 VPWR \$238 VGND \$214 VPWR \$215 VGND sky130_fd_sc_hd__nor2_1
X$760 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$761 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$762 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$763 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$764 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$765 VPWR \$232 VPWR VGND \$239 \$225 VGND sky130_fd_sc_hd__nand2_1
X$766 VPWR VGND \$218 VPWR \$198 \$217 \$239 VGND sky130_fd_sc_hd__a21o_1
X$767 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$768 VPWR \$225 VPWR VGND \$217 \$218 \$198 VGND sky130_fd_sc_hd__nand3_1
X$769 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$770 VGND \$35 \$240 \$168 \$232 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$771 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$772 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$773 VGND \$187 \$190 \$208 \$198 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$774 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$775 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$776 VGND \$35 \$196 \$188 \$191 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$777 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$778 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$779 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$780 VPWR VGND \$240 \$217 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$781 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$782 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$783 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$784 VPWR sel2[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$785 VPWR \$192 VGND VPWR sel2[0] VGND sky130_fd_sc_hd__clkbuf_1
X$786 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$787 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$788 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$789 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$790 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$791 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$792 VPWR \$132 VGND VPWR \$126 VGND sky130_fd_sc_hd__clkbuf_1
X$793 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$794 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$795 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$796 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$797 VPWR \$85 VGND \$44 VPWR \$96 VGND sky130_fd_sc_hd__nor2_1
X$798 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$799 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$800 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$801 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$802 VPWR \$64 VGND VPWR \$97 VGND sky130_fd_sc_hd__dlygate4sd1_1
X$803 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$804 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$805 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$806 VGND \$100 \$128 \$108 \$32 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$807 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$808 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$809 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$810 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$811 VGND \$35 \$119 \$60 \$131 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$812 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$813 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$814 VPWR \$134 VPWR \$112 VGND \$119 VGND sky130_fd_sc_hd__xnor2_1
X$815 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$816 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$817 VPWR VGND VPWR \$39 \$120 VGND sky130_fd_sc_hd__inv_4
X$818 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$819 VPWR \$124 VGND \$121 VPWR \$128 VGND sky130_fd_sc_hd__nor2_1
X$820 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$821 VGND \$121 \$39 \$128 VPWR VPWR VGND sky130_fd_sc_hd__dfxtp_1
X$822 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$823 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$824 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$825 VGND \$35 \$38 \$138 \$125 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_4
X$826 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$827 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$828 VPWR sel[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$829 VPWR \$135 VGND VPWR sel[1] VGND sky130_fd_sc_hd__clkbuf_1
X$830 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$831 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$832 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$833 VGND \$35 \$140 \$60 \$132 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_2
X$834 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$835 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$836 VGND \$136 \$142 \$144 \$106 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$837 VGND \$126 \$140 \$133 \$106 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$838 VPWR \$127 \$140 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$839 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$840 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$841 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$842 VPWR \$140 \$145 VGND \$142 VPWR \$38 VGND sky130_fd_sc_hd__nor3_1
X$843 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$844 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$845 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$846 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$847 VPWR \$146 VGND \$142 VPWR \$143 VGND sky130_fd_sc_hd__nor2_1
X$848 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$849 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$850 VPWR VGND \$109 \$137 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$851 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$852 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$853 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$854 VGND \$137 \$141 \$138 \$80 \$134 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2ai_2
X$855 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$856 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$857 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$858 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$859 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$860 VGND \$35 \$147 \$138 \$139 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_1
X$861 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$862 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$863 VPWR VGND \$128 VPWR \$54 VGND sky130_fd_sc_hd__buf_2
X$864 VGND \$35 \$152 \$138 \$135 VPWR VPWR VGND sky130_fd_sc_hd__dfstp_1
X$865 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$866 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$867 VPWR \$35 VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$868 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$869 VPWR VGND \$43 \$160 VPWR VGND sky130_fd_sc_hd__clkinv_4
X$870 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$871 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
.ENDS caravel_clocking

.SUBCKT sky130_fd_sc_hd__dlymetal6s2s_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__dlymetal6s2s_1

.SUBCKT sky130_fd_sc_hd__clkbuf_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_4

.SUBCKT sky130_fd_sc_hd__dfstp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_2

.SUBCKT sky130_fd_sc_hd__nor3b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3b_1

.SUBCKT sky130_fd_sc_hd__o211a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211a_1

.SUBCKT sky130_fd_sc_hd__dfrtp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_2

.SUBCKT sky130_fd_sc_hd__or2b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2b_1

.SUBCKT sky130_fd_sc_hd__nand2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__buf_12 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_12

.SUBCKT sky130_fd_sc_hd__a21bo_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21bo_1

.SUBCKT sky130_fd_sc_hd__buf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__mux2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_2

.SUBCKT sky130_fd_sc_hd__o211ai_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211ai_4

.SUBCKT sky130_fd_sc_hd__nor3b_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3b_2

.SUBCKT sky130_fd_sc_hd__and2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__and2_1

.SUBCKT sky130_fd_sc_hd__conb_1 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__buf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__inv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__o21bai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21bai_1

.SUBCKT sky130_fd_sc_hd__nand3b_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nand3b_1

.SUBCKT sky130_fd_sc_hd__clkdlybuf4s25_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkdlybuf4s25_1

.SUBCKT sky130_fd_sc_hd__dfstp_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_4

.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o2bb2ai_2

.SUBCKT sky130_fd_sc_hd__a21o_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21o_1

.SUBCKT sky130_fd_sc_hd__clkinv_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_4

.SUBCKT sky130_fd_sc_hd__o21a_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21a_1

.SUBCKT sky130_fd_sc_hd__nand2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_1

.SUBCKT sky130_fd_sc_hd__dfrtp_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_4

.SUBCKT sky130_fd_sc_hd__nor3_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nor3_1

.SUBCKT sky130_fd_sc_hd__clkbuf_16 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_16

.SUBCKT sky130_fd_sc_hd__dfrtn_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtn_1

.SUBCKT sky130_fd_sc_hd__inv_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_4

.SUBCKT sky130_fd_sc_hd__xor2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__xor2_1

.SUBCKT sky130_fd_sc_hd__decap_12 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__dfrtp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_1

.SUBCKT sky130_fd_sc_hd__nor2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_1

.SUBCKT sky130_fd_sc_hd__diode_2 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__dfxtp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__dfxtp_1

.SUBCKT sky130_fd_sc_hd__nand3_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__nand3_1

.SUBCKT sky130_fd_sc_hd__clkbuf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__fill_2 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__mux2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 nc_1 nc_2
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__xnor2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__xnor2_1

.SUBCKT sky130_fd_sc_hd__clkbuf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__decap_8 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__fill_1 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__dfstp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfstp_1

.SUBCKT sky130_fd_sc_hd__decap_6 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__decap_4 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__o21ai_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ai_1

.SUBCKT sky130_fd_sc_hd__dlygate4sd1_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__dlygate4sd1_1

.SUBCKT sky130_fd_sc_hd__decap_3 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__clkinv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_2
