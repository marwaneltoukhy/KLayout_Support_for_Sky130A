*SPICE netlist created from verilog structural netlist module gpio_defaults_block by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /home/marwan/klayout_lvs/lvs/test_cases/gpio_defaults_block/sky130_fd_sc_hd.spice

.subckt gpio_defaults_block VGND VPWR gpio_defaults[0] gpio_defaults[1] gpio_defaults[2] gpio_defaults[3] gpio_defaults[4]
+ gpio_defaults[5] gpio_defaults[6] gpio_defaults[7] gpio_defaults[8] gpio_defaults[9] gpio_defaults[10] gpio_defaults[11] gpio_defaults[12]
+ 

XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_10 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_6 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_7 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X\gpio_default_value[0]  VGND VGND VPWR VPWR \gpio_defaults_high[0]\ \gpio_defaults_low[0]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[10]  VGND VGND VPWR VPWR \gpio_defaults_high[10]\ \gpio_defaults_low[10]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[11]  VGND VGND VPWR VPWR \gpio_defaults_high[11]\ \gpio_defaults_low[11]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[12]  VGND VGND VPWR VPWR \gpio_defaults_high[12]\ \gpio_defaults_low[12]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[1]  VGND VGND VPWR VPWR \gpio_defaults_high[1]\ \gpio_defaults_low[1]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[2]  VGND VGND VPWR VPWR \gpio_defaults_high[2]\ \gpio_defaults_low[2]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[3]  VGND VGND VPWR VPWR \gpio_defaults_high[3]\ \gpio_defaults_low[3]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[4]  VGND VGND VPWR VPWR \gpio_defaults_high[4]\ \gpio_defaults_low[4]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[5]  VGND VGND VPWR VPWR \gpio_defaults_high[5]\ \gpio_defaults_low[5]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[6]  VGND VGND VPWR VPWR \gpio_defaults_high[6]\ \gpio_defaults_low[6]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[7]  VGND VGND VPWR VPWR \gpio_defaults_high[7]\ \gpio_defaults_low[7]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[8]  VGND VGND VPWR VPWR \gpio_defaults_high[8]\ \gpio_defaults_low[8]\ sky130_fd_sc_hd__conb_1
X\gpio_default_value[9]  VGND VGND VPWR VPWR \gpio_defaults_high[9]\ \gpio_defaults_low[9]\ sky130_fd_sc_hd__conb_1

.ends
.end
