*SPICE netlist created from verilog structural netlist module housekeeping by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /home/marwan/klayout_lvs/lvs/test_cases/housekeeping/sky130_fd_sc_hd.spice

.subckt housekeeping VGND VPWR debug_in debug_mode debug_oeb debug_out pad_flash_clk
+ pad_flash_clk_oeb pad_flash_csb pad_flash_csb_oeb pad_flash_io0_di pad_flash_io0_do pad_flash_io0_ieb pad_flash_io0_oeb pad_flash_io1_di
+ pad_flash_io1_do pad_flash_io1_ieb pad_flash_io1_oeb pll_bypass pll_dco_ena pll_ena porb qspi_enabled
+ reset ser_rx ser_tx serial_clock serial_data_1 serial_data_2 serial_load serial_resetn
+ spi_csb spi_enabled spi_sck spi_sdi spi_sdo spi_sdoenb spimemio_flash_clk spimemio_flash_csb
+ spimemio_flash_io0_di spimemio_flash_io0_do spimemio_flash_io0_oeb spimemio_flash_io1_di spimemio_flash_io1_do spimemio_flash_io1_oeb spimemio_flash_io2_di spimemio_flash_io2_do
+ spimemio_flash_io2_oeb spimemio_flash_io3_di spimemio_flash_io3_do spimemio_flash_io3_oeb sram_ro_clk sram_ro_csb trap uart_enabled
+ user_clock usr1_vcc_pwrgood usr1_vdd_pwrgood usr2_vcc_pwrgood usr2_vdd_pwrgood wb_ack_o wb_clk_i wb_cyc_i
+ wb_rstn_i wb_stb_i wb_we_i irq[0] irq[1] irq[2] mask_rev_in[0] mask_rev_in[1]
+ mask_rev_in[2] mask_rev_in[3] mask_rev_in[4] mask_rev_in[5] mask_rev_in[6] mask_rev_in[7] mask_rev_in[8] mask_rev_in[9]
+ mask_rev_in[10] mask_rev_in[11] mask_rev_in[12] mask_rev_in[13] mask_rev_in[14] mask_rev_in[15] mask_rev_in[16] mask_rev_in[17]
+ mask_rev_in[18] mask_rev_in[19] mask_rev_in[20] mask_rev_in[21] mask_rev_in[22] mask_rev_in[23] mask_rev_in[24] mask_rev_in[25]
+ mask_rev_in[26] mask_rev_in[27] mask_rev_in[28] mask_rev_in[29] mask_rev_in[30] mask_rev_in[31] mgmt_gpio_in[0] mgmt_gpio_in[1]
+ mgmt_gpio_in[2] mgmt_gpio_in[3] mgmt_gpio_in[4] mgmt_gpio_in[5] mgmt_gpio_in[6] mgmt_gpio_in[7] mgmt_gpio_in[8] mgmt_gpio_in[9]
+ mgmt_gpio_in[10] mgmt_gpio_in[11] mgmt_gpio_in[12] mgmt_gpio_in[13] mgmt_gpio_in[14] mgmt_gpio_in[15] mgmt_gpio_in[16] mgmt_gpio_in[17]
+ mgmt_gpio_in[18] mgmt_gpio_in[19] mgmt_gpio_in[20] mgmt_gpio_in[21] mgmt_gpio_in[22] mgmt_gpio_in[23] mgmt_gpio_in[24] mgmt_gpio_in[25]
+ mgmt_gpio_in[26] mgmt_gpio_in[27] mgmt_gpio_in[28] mgmt_gpio_in[29] mgmt_gpio_in[30] mgmt_gpio_in[31] mgmt_gpio_in[32] mgmt_gpio_in[33]
+ mgmt_gpio_in[34] mgmt_gpio_in[35] mgmt_gpio_in[36] mgmt_gpio_in[37] mgmt_gpio_oeb[0] mgmt_gpio_oeb[1] mgmt_gpio_oeb[2] mgmt_gpio_oeb[3]
+ mgmt_gpio_oeb[4] mgmt_gpio_oeb[5] mgmt_gpio_oeb[6] mgmt_gpio_oeb[7] mgmt_gpio_oeb[8] mgmt_gpio_oeb[9] mgmt_gpio_oeb[10] mgmt_gpio_oeb[11]
+ mgmt_gpio_oeb[12] mgmt_gpio_oeb[13] mgmt_gpio_oeb[14] mgmt_gpio_oeb[15] mgmt_gpio_oeb[16] mgmt_gpio_oeb[17] mgmt_gpio_oeb[18] mgmt_gpio_oeb[19]
+ mgmt_gpio_oeb[20] mgmt_gpio_oeb[21] mgmt_gpio_oeb[22] mgmt_gpio_oeb[23] mgmt_gpio_oeb[24] mgmt_gpio_oeb[25] mgmt_gpio_oeb[26] mgmt_gpio_oeb[27]
+ mgmt_gpio_oeb[28] mgmt_gpio_oeb[29] mgmt_gpio_oeb[30] mgmt_gpio_oeb[31] mgmt_gpio_oeb[32] mgmt_gpio_oeb[33] mgmt_gpio_oeb[34] mgmt_gpio_oeb[35]
+ mgmt_gpio_oeb[36] mgmt_gpio_oeb[37] mgmt_gpio_out[0] mgmt_gpio_out[1] mgmt_gpio_out[2] mgmt_gpio_out[3] mgmt_gpio_out[4] mgmt_gpio_out[5]
+ mgmt_gpio_out[6] mgmt_gpio_out[7] mgmt_gpio_out[8] mgmt_gpio_out[9] mgmt_gpio_out[10] mgmt_gpio_out[11] mgmt_gpio_out[12] mgmt_gpio_out[13]
+ mgmt_gpio_out[14] mgmt_gpio_out[15] mgmt_gpio_out[16] mgmt_gpio_out[17] mgmt_gpio_out[18] mgmt_gpio_out[19] mgmt_gpio_out[20] mgmt_gpio_out[21]
+ mgmt_gpio_out[22] mgmt_gpio_out[23] mgmt_gpio_out[24] mgmt_gpio_out[25] mgmt_gpio_out[26] mgmt_gpio_out[27] mgmt_gpio_out[28] mgmt_gpio_out[29]
+ mgmt_gpio_out[30] mgmt_gpio_out[31] mgmt_gpio_out[32] mgmt_gpio_out[33] mgmt_gpio_out[34] mgmt_gpio_out[35] mgmt_gpio_out[36] mgmt_gpio_out[37]
+ pll90_sel[0] pll90_sel[1] pll90_sel[2] pll_div[0] pll_div[1] pll_div[2] pll_div[3] pll_div[4]
+ pll_sel[0] pll_sel[1] pll_sel[2] pll_trim[0] pll_trim[1] pll_trim[2] pll_trim[3] pll_trim[4]
+ pll_trim[5] pll_trim[6] pll_trim[7] pll_trim[8] pll_trim[9] pll_trim[10] pll_trim[11] pll_trim[12]
+ pll_trim[13] pll_trim[14] pll_trim[15] pll_trim[16] pll_trim[17] pll_trim[18] pll_trim[19] pll_trim[20]
+ pll_trim[21] pll_trim[22] pll_trim[23] pll_trim[24] pll_trim[25] pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2]
+ pwr_ctrl_out[3] sram_ro_addr[0] sram_ro_addr[1] sram_ro_addr[2] sram_ro_addr[3] sram_ro_addr[4] sram_ro_addr[5] sram_ro_addr[6]
+ sram_ro_addr[7] sram_ro_data[0] sram_ro_data[1] sram_ro_data[2] sram_ro_data[3] sram_ro_data[4] sram_ro_data[5] sram_ro_data[6]
+ sram_ro_data[7] sram_ro_data[8] sram_ro_data[9] sram_ro_data[10] sram_ro_data[11] sram_ro_data[12] sram_ro_data[13] sram_ro_data[14]
+ sram_ro_data[15] sram_ro_data[16] sram_ro_data[17] sram_ro_data[18] sram_ro_data[19] sram_ro_data[20] sram_ro_data[21] sram_ro_data[22]
+ sram_ro_data[23] sram_ro_data[24] sram_ro_data[25] sram_ro_data[26] sram_ro_data[27] sram_ro_data[28] sram_ro_data[29] sram_ro_data[30]
+ sram_ro_data[31] wb_adr_i[0] wb_adr_i[1] wb_adr_i[2] wb_adr_i[3] wb_adr_i[4] wb_adr_i[5] wb_adr_i[6]
+ wb_adr_i[7] wb_adr_i[8] wb_adr_i[9] wb_adr_i[10] wb_adr_i[11] wb_adr_i[12] wb_adr_i[13] wb_adr_i[14]
+ wb_adr_i[15] wb_adr_i[16] wb_adr_i[17] wb_adr_i[18] wb_adr_i[19] wb_adr_i[20] wb_adr_i[21] wb_adr_i[22]
+ wb_adr_i[23] wb_adr_i[24] wb_adr_i[25] wb_adr_i[26] wb_adr_i[27] wb_adr_i[28] wb_adr_i[29] wb_adr_i[30]
+ wb_adr_i[31] wb_dat_i[0] wb_dat_i[1] wb_dat_i[2] wb_dat_i[3] wb_dat_i[4] wb_dat_i[5] wb_dat_i[6]
+ wb_dat_i[7] wb_dat_i[8] wb_dat_i[9] wb_dat_i[10] wb_dat_i[11] wb_dat_i[12] wb_dat_i[13] wb_dat_i[14]
+ wb_dat_i[15] wb_dat_i[16] wb_dat_i[17] wb_dat_i[18] wb_dat_i[19] wb_dat_i[20] wb_dat_i[21] wb_dat_i[22]
+ wb_dat_i[23] wb_dat_i[24] wb_dat_i[25] wb_dat_i[26] wb_dat_i[27] wb_dat_i[28] wb_dat_i[29] wb_dat_i[30]
+ wb_dat_i[31] wb_dat_o[0] wb_dat_o[1] wb_dat_o[2] wb_dat_o[3] wb_dat_o[4] wb_dat_o[5] wb_dat_o[6]
+ wb_dat_o[7] wb_dat_o[8] wb_dat_o[9] wb_dat_o[10] wb_dat_o[11] wb_dat_o[12] wb_dat_o[13] wb_dat_o[14]
+ wb_dat_o[15] wb_dat_o[16] wb_dat_o[17] wb_dat_o[18] wb_dat_o[19] wb_dat_o[20] wb_dat_o[21] wb_dat_o[22]
+ wb_dat_o[23] wb_dat_o[24] wb_dat_o[25] wb_dat_o[26] wb_dat_o[27] wb_dat_o[28] wb_dat_o[29] wb_dat_o[30]
+ wb_dat_o[31] wb_sel_i[0] wb_sel_i[1] wb_sel_i[2] wb_sel_i[3] 

XANTENNA_0 user_clock VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_1 wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_10 _0113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_100 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_101 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_102 net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_103 net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_104 net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_105 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_106 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_107 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_108 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_109 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 _0115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_110 net77 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_111 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_112 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_113 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_114 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_115 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_116 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_117 net85 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_118 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_119 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 _0115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_120 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_121 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_122 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_123 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_124 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_125 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_126 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_127 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_128 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_129 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_13 _0115_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_130 net87 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_131 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_132 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_133 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_134 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_135 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_136 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_137 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_138 _0085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_139 _0093_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 _0117_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_140 _0107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_141 _0107_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_142 _0109_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_143 _0134_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_144 _0144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_145 _0144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_146 _0144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_147 _0152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_148 _0152_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_149 _1023_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_15 _0119_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_150 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_151 _1106_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_152 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_153 _1181_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_154 _1245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_155 _1245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_156 _1245_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_157 _1275_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_158 _1292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_159 _1292_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_16 _0121_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_160 _1293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_161 _2032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_162 _2045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_163 _2045_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_164 _2239_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_165 _2306_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_166 _2338_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_167 _2542_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_168 _2554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_169 _2554_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_17 _0123_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_170 _2637_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_171 _2664_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_172 _3010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_173 _3010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_174 _3435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_175 _3600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_176 _4268_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_177 _4421_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_178 _4423_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_179 \gpio_configure[19][6]\ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_18 _0125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_180 \hkspi.idata[2]\ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_181 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_182 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_183 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_184 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_185 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_186 net201 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_187 net205 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_188 net206 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_189 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_19 _0130_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_190 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_191 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_192 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_193 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_194 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_195 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_196 net313 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_197 net78 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_198 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_199 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_2 _0079_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_20 _0132_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_200 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_201 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_202 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_203 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_204 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_205 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_206 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_207 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_208 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_209 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 _0142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_210 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_211 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_212 _1235_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_213 _1861_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_214 _2414_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_215 _2416_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_216 _4410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_217 net368 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_218 net307 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_22 _0142_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 _0148_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_24 _0150_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_25 _1043_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_26 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_27 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_28 _1047_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_29 _1158_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_3 _0083_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_30 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_31 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_32 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_33 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_34 _1256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_35 _1267_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_36 _1283_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_37 _1311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_38 _1313_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_39 _1320_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_4 _0103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_40 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_41 _1329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_42 _1329_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_43 _1336_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_44 _1345_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_45 _1367_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_46 _1387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_47 _1399_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_48 _1411_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_49 _1870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _0103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_50 _1890_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_51 _1895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_52 _1899_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_53 _1905_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_54 _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_55 _1988_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_56 _1993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_57 _2033_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_58 _2037_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_59 _2052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_6 _0103_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_60 _2060_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_61 _2072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_62 _2072_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_63 _2075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_64 _2224_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_65 _2342_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_66 _2413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_67 _2417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_68 _2440_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_69 _2443_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_7 _0105_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_70 _2464_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_71 _2484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_72 _2520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_73 _2520_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_74 _2563_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_75 _2567_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_76 _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_77 _2593_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_78 _2645_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_79 _2816_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_8 _0111_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_80 _2977_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_81 _2998_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_82 _3151_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_83 _3309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_84 _4000_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_85 _4206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_86 _4206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_87 _4417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_88 _4432_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_89 _4436_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_9 _0113_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_90 clknet_3_6_0_wb_clk_i VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_91 \hkspi.idata[5]\ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_92 \mgmt_gpio_data[9]\ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_93 net207 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_94 net245 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_95 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_96 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_97 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_98 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_99 net312 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_112_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_161_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_161_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_162_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_162_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_177_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_185_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_187_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4443_ \mgmt_gpio_data[32]\ net80 net79 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[32]\ sky130_fd_sc_hd__mux2_1
X_4444_ \mgmt_gpio_data[33]\ net78 net79 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[33]\ sky130_fd_sc_hd__mux2_1
X_4445_ \mgmt_gpio_data[10]\ net58 \hkspi.pass_thru_user\ VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[10]\ sky130_fd_sc_hd__mux2_1
X_4446_ \mgmt_gpio_data[9]\ clknet_2_3_0_mgmt_gpio_in[4] \hkspi.pass_thru_user\ VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[9]\ sky130_fd_sc_hd__mux2_1
X_4447_ \mgmt_gpio_data[8]\ net67 \hkspi.pass_thru_user_delay\ VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[8]\ sky130_fd_sc_hd__mux2_1
X_4448_ \mgmt_gpio_data[6]\ net77 net126 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[6]\ sky130_fd_sc_hd__mux2_1
X_4449_ \mgmt_gpio_data[15]\ user_clock clk2_output_dest VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[15]\ sky130_fd_sc_hd__mux2_1
X_4450_ \mgmt_gpio_data[14]\ clknet_3_6_0_wb_clk_i clk1_output_dest VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[14]\ sky130_fd_sc_hd__mux2_1
X_4451_ \mgmt_gpio_data[13]\ net125 trap_output_dest VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_out_pre[13]\ sky130_fd_sc_hd__mux2_1
X_4452_ _0063_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__clkinv_2
X_4453_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__buf_12
X_4454_ _1022_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__buf_12
X_4455_ _0073_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__inv_2
X_4456_ wbbd_busy VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__inv_2
X_4457_ _1025_ _0078_ _0077_ VGND VGND VPWR 
+ VPWR
+ _1026_ sky130_fd_sc_hd__a21o_1
X_4458_ _1024_ _0075_ _1026_ VGND VGND VPWR 
+ VPWR
+ _1027_ sky130_fd_sc_hd__or3_1
X_4459_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__clkbuf_8
X_4460_ _0067_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__clkinv_2
X_4461_ _0065_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__clkinv_2
X_4462_ _1029_ _1030_ _0071_ _0069_ VGND VGND 
+ VPWR
+ VPWR _1031_ sky130_fd_sc_hd__or4_4
X_4463_ _1028_ _1031_ VGND VGND VPWR VPWR 
+ _1032_
+ sky130_fd_sc_hd__or2_4
X_4464_ _1023_ _1032_ VGND VGND VPWR VPWR 
+ _1033_
+ sky130_fd_sc_hd__or2_1
X_4465_ _1033_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__buf_2
X_4466_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__clkinv_2
X_4467_ serial_bb_data_2 _1034_ \cdata[6]\ _1035_ VGND VGND 
+ VPWR
+ VPWR _1019_ sky130_fd_sc_hd__a22o_1
X_4468_ _0075_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__inv_2
X_4469_ _1025_ _0078_ _0077_ VGND VGND VPWR 
+ VPWR
+ _1037_ sky130_fd_sc_hd__a21bo_1
X_4470_ _0073_ _1036_ _1037_ VGND VGND VPWR 
+ VPWR
+ _1038_ sky130_fd_sc_hd__or3_1
X_4471_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__buf_8
X_4472_ _0071_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__clkinv_2
X_4473_ _0069_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__clkinv_2
X_4474_ _1029_ _1030_ _1040_ _1041_ VGND VGND 
+ VPWR
+ VPWR _1042_ sky130_fd_sc_hd__or4_4
X_4475_ _1022_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__buf_12
X_4476_ _1039_ _1042_ _1043_ VGND VGND VPWR 
+ VPWR
+ _1044_ sky130_fd_sc_hd__or3_1
X_4477_ \cdata[0]\ hkspi_disable _1044_ VGND VGND VPWR 
+ VPWR
+ _1045_ sky130_fd_sc_hd__mux2_1
X_4478_ _1045_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__clkbuf_1
X_4479_ _1029_ _1030_ _1040_ _0069_ VGND VGND 
+ VPWR
+ VPWR _1046_ sky130_fd_sc_hd__or4_4
X_4480_ _1028_ _1046_ VGND VGND VPWR VPWR 
+ _1047_
+ sky130_fd_sc_hd__or2_4
X_4481_ _1043_ _1047_ VGND VGND VPWR VPWR 
+ _1048_
+ sky130_fd_sc_hd__or2_2
X_4482_ net364 clk1_output_dest _1048_ VGND VGND VPWR 
+ VPWR
+ _1049_ sky130_fd_sc_hd__mux2_1
X_4483_ _1049_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__clkbuf_1
X_4484_ serial_bb_enable _1034_ net366 _1035_ VGND VGND 
+ VPWR
+ VPWR _1016_ sky130_fd_sc_hd__a22o_1
X_4485_ \cdata[1]\ clk2_output_dest _1048_ VGND VGND VPWR 
+ VPWR
+ _1050_ sky130_fd_sc_hd__mux2_1
X_4486_ _1050_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__clkbuf_1
X_4487_ _1024_ _0075_ _1037_ VGND VGND VPWR 
+ VPWR
+ _1051_ sky130_fd_sc_hd__or3_1
X_4488_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__buf_6
X_4489_ _0071_ _0069_ _0067_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1053_ sky130_fd_sc_hd__or4_4
X_4490_ _1052_ _1053_ VGND VGND VPWR VPWR 
+ _1054_
+ sky130_fd_sc_hd__or2_4
X_4491_ _1023_ _1054_ VGND VGND VPWR VPWR 
+ _1055_
+ sky130_fd_sc_hd__or2_1
X_4492_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__buf_2
X_4493_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__inv_2
X_4494_ \gpio_configure[25][7]\ _1056_ \cdata[7]\ _1057_ VGND VGND 
+ VPWR
+ VPWR _1014_ sky130_fd_sc_hd__a22o_1
X_4495_ \gpio_configure[25][6]\ _1056_ \cdata[6]\ _1057_ VGND VGND 
+ VPWR
+ VPWR _1013_ sky130_fd_sc_hd__a22o_1
X_4496_ \gpio_configure[25][5]\ _1056_ \cdata[5]\ _1057_ VGND VGND 
+ VPWR
+ VPWR _1012_ sky130_fd_sc_hd__a22o_1
X_4497_ \gpio_configure[25][4]\ _1056_ net359 _1057_ VGND VGND 
+ VPWR
+ VPWR _1011_ sky130_fd_sc_hd__a22o_1
X_4498_ \gpio_configure[25][3]\ _1056_ net361 _1057_ VGND VGND 
+ VPWR
+ VPWR _1010_ sky130_fd_sc_hd__a22o_1
X_4499_ \gpio_configure[25][2]\ _1056_ net363 _1057_ VGND VGND 
+ VPWR
+ VPWR _1009_ sky130_fd_sc_hd__a22o_1
X_4500_ \gpio_configure[25][1]\ _1056_ net366 _1057_ VGND VGND 
+ VPWR
+ VPWR _1008_ sky130_fd_sc_hd__a22o_1
X_4501_ \gpio_configure[25][0]\ _1056_ net367 _1057_ VGND VGND 
+ VPWR
+ VPWR _1007_ sky130_fd_sc_hd__a22o_1
X_4502_ _0071_ _0069_ _0067_ _1030_ VGND VGND 
+ VPWR
+ VPWR _1058_ sky130_fd_sc_hd__or4_4
X_4503_ _1052_ _1058_ VGND VGND VPWR VPWR 
+ _1059_
+ sky130_fd_sc_hd__or2_4
X_4504_ _1043_ _1059_ VGND VGND VPWR VPWR 
+ _1060_
+ sky130_fd_sc_hd__or2_1
X_4505_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__clkbuf_2
X_4506_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__inv_2
X_4507_ \gpio_configure[26][12]\ _1061_ net359 _1062_ VGND VGND 
+ VPWR
+ VPWR _1006_ sky130_fd_sc_hd__a22o_1
X_4508_ \gpio_configure[26][11]\ _1061_ net361 _1062_ VGND VGND 
+ VPWR
+ VPWR _1005_ sky130_fd_sc_hd__a22o_1
X_4509_ \gpio_configure[26][10]\ _1061_ net363 _1062_ VGND VGND 
+ VPWR
+ VPWR _1004_ sky130_fd_sc_hd__a22o_1
X_4510_ \gpio_configure[26][9]\ _1061_ net365 _1062_ VGND VGND 
+ VPWR
+ VPWR _1003_ sky130_fd_sc_hd__a22o_1
X_4511_ \gpio_configure[26][8]\ _1061_ net367 _1062_ VGND VGND 
+ VPWR
+ VPWR _1002_ sky130_fd_sc_hd__a22o_1
X_4512_ serial_bb_clock _1034_ net359 _1035_ VGND VGND 
+ VPWR
+ VPWR _1001_ sky130_fd_sc_hd__a22o_2
X_4513_ _1040_ _0069_ _1029_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1063_ sky130_fd_sc_hd__or4_4
X_4514_ _0073_ _0075_ _1026_ VGND VGND VPWR 
+ VPWR
+ _1064_ sky130_fd_sc_hd__or3_1
X_4515_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__buf_8
X_4516_ _1063_ _1065_ VGND VGND VPWR VPWR 
+ _1066_
+ sky130_fd_sc_hd__or2_2
X_4517_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__inv_2
X_4518_ net204 _1067_ net367 _1066_ _0063_ VGND 
+ VGND
+ VPWR VPWR _1000_ sky130_fd_sc_hd__o221a_1
X_4519_ _1046_ _1065_ _1043_ VGND VGND VPWR 
+ VPWR
+ _1068_ sky130_fd_sc_hd__or3_1
X_4520_ net367 reset_reg _1068_ VGND VGND VPWR 
+ VPWR
+ _1069_ sky130_fd_sc_hd__mux2_1
X_4521_ _1069_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__clkbuf_1
X_4522_ _0067_ _1030_ _0071_ _1041_ VGND VGND 
+ VPWR
+ VPWR _1070_ sky130_fd_sc_hd__or4_4
X_4523_ _1028_ _1070_ VGND VGND VPWR VPWR 
+ _1071_
+ sky130_fd_sc_hd__or2_4
X_4524_ _1023_ _1071_ VGND VGND VPWR VPWR 
+ _1072_
+ sky130_fd_sc_hd__or2_1
X_4525_ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__clkbuf_4
X_4526_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__inv_2
X_4527_ net323 _1073_ \cdata[7]\ _1074_ VGND VGND 
+ VPWR
+ VPWR _0998_ sky130_fd_sc_hd__a22o_1
X_4528_ net322 _1073_ \cdata[6]\ _1074_ VGND VGND 
+ VPWR
+ VPWR _0997_ sky130_fd_sc_hd__a22o_1
X_4529_ net321 _1073_ \cdata[5]\ _1074_ VGND VGND 
+ VPWR
+ VPWR _0996_ sky130_fd_sc_hd__a22o_1
X_4530_ net320 _1073_ net359 _1074_ VGND VGND 
+ VPWR
+ VPWR _0995_ sky130_fd_sc_hd__a22o_1
X_4531_ net319 _1073_ net361 _1074_ VGND VGND 
+ VPWR
+ VPWR _0994_ sky130_fd_sc_hd__a22o_1
X_4532_ net318 _1073_ net363 _1074_ VGND VGND 
+ VPWR
+ VPWR _0993_ sky130_fd_sc_hd__a22o_1
X_4533_ net317 _1073_ net365 _1074_ VGND VGND 
+ VPWR
+ VPWR _0992_ sky130_fd_sc_hd__a22o_1
X_4534_ net316 _1073_ net367 _1074_ VGND VGND 
+ VPWR
+ VPWR _0991_ sky130_fd_sc_hd__a22o_1
X_4535_ _0067_ _0065_ _0071_ _1041_ VGND VGND 
+ VPWR
+ VPWR _1075_ sky130_fd_sc_hd__or4_4
X_4536_ _1028_ _1075_ VGND VGND VPWR VPWR 
+ _1076_
+ sky130_fd_sc_hd__or2_2
X_4537_ _1043_ _1076_ VGND VGND VPWR VPWR 
+ _1077_
+ sky130_fd_sc_hd__or2_2
X_4538_ net367 net325 _1077_ VGND VGND VPWR 
+ VPWR
+ _1078_ sky130_fd_sc_hd__mux2_1
X_4539_ _1078_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__clkbuf_1
X_4540_ net365 net324 _1077_ VGND VGND VPWR 
+ VPWR
+ _1079_ sky130_fd_sc_hd__mux2_1
X_4541_ _1079_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__clkbuf_1
X_4542_ \wbbd_state[6]\ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__clkinv_2
X_4543_ \wbbd_state[5]\ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__inv_2
X_4544_ \wbbd_state[7]\ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__inv_2
X_4545_ \wbbd_state[8]\ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__inv_2
X_4546_ \wbbd_state[9]\ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__inv_2
X_4547_ _1082_ _1083_ _1084_ VGND VGND VPWR 
+ VPWR
+ _1085_ sky130_fd_sc_hd__and3_1
X_4548_ _1085_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__buf_12
X_4549_ _1081_ _0169_ VGND VGND VPWR VPWR 
+ _1086_
+ sky130_fd_sc_hd__nand2_8
X_4550_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__inv_6
X_4551_ \wbbd_state[6]\ _1086_ VGND VGND VPWR VPWR 
+ _1088_
+ sky130_fd_sc_hd__or2_1
X_4552_ _1080_ _1087_ wbbd_write _4442_ _1088_ VGND 
+ VGND
+ VPWR VPWR _0988_ sky130_fd_sc_hd__a32o_1
X_4553_ _1040_ _0069_ _0067_ _1030_ VGND VGND 
+ VPWR
+ VPWR _1089_ sky130_fd_sc_hd__or4_4
X_4554_ _1065_ _1089_ _1043_ VGND VGND VPWR 
+ VPWR
+ _1090_ sky130_fd_sc_hd__or3_1
X_4555_ net367 net263 _1090_ VGND VGND VPWR 
+ VPWR
+ _1091_ sky130_fd_sc_hd__mux2_1
X_4556_ _1091_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__clkbuf_1
X_4557_ _1028_ _1053_ VGND VGND VPWR VPWR 
+ _1092_
+ sky130_fd_sc_hd__or2_2
X_4558_ _1043_ _1092_ VGND VGND VPWR VPWR 
+ _1093_
+ sky130_fd_sc_hd__or2_1
X_4559_ net365 net291 _1093_ VGND VGND VPWR 
+ VPWR
+ _1094_ sky130_fd_sc_hd__mux2_1
X_4560_ _1094_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__clkbuf_1
X_4561_ net367 net290 _1093_ VGND VGND VPWR 
+ VPWR
+ _1095_ sky130_fd_sc_hd__mux2_1
X_4562_ _1095_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_1
X_4563_ _1042_ _1065_ VGND VGND VPWR VPWR 
+ _1096_
+ sky130_fd_sc_hd__or2_4
X_4564_ _1023_ _1096_ VGND VGND VPWR VPWR 
+ _1097_
+ sky130_fd_sc_hd__or2_1
X_4565_ _1097_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__buf_2
X_4566_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__clkinv_2
X_4567_ net289 _1098_ \cdata[7]\ _1099_ VGND VGND 
+ VPWR
+ VPWR _0984_ sky130_fd_sc_hd__a22o_1
X_4568_ net288 _1098_ \cdata[6]\ _1099_ VGND VGND 
+ VPWR
+ VPWR _0983_ sky130_fd_sc_hd__a22o_1
X_4569_ net287 _1098_ \cdata[5]\ _1099_ VGND VGND 
+ VPWR
+ VPWR _0982_ sky130_fd_sc_hd__a22o_1
X_4570_ net286 _1098_ net359 _1099_ VGND VGND 
+ VPWR
+ VPWR _0981_ sky130_fd_sc_hd__a22o_1
X_4571_ net284 _1098_ net361 _1099_ VGND VGND 
+ VPWR
+ VPWR _0980_ sky130_fd_sc_hd__a22o_1
X_4572_ net283 _1098_ net363 _1099_ VGND VGND 
+ VPWR
+ VPWR _0979_ sky130_fd_sc_hd__a22o_1
X_4573_ net282 _1098_ net365 _1099_ VGND VGND 
+ VPWR
+ VPWR _0978_ sky130_fd_sc_hd__a22o_1
X_4574_ net281 _1098_ net367 _1099_ VGND VGND 
+ VPWR
+ VPWR _0977_ sky130_fd_sc_hd__a22o_1
X_4575_ _1040_ _1041_ _1029_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1100_ sky130_fd_sc_hd__or4_4
X_4576_ _1065_ _1100_ VGND VGND VPWR VPWR 
+ _1101_
+ sky130_fd_sc_hd__or2_4
X_4577_ _1023_ _1101_ VGND VGND VPWR VPWR 
+ _1102_
+ sky130_fd_sc_hd__or2_1
X_4578_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__clkbuf_4
X_4579_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__clkinv_2
X_4580_ net280 _1103_ \cdata[7]\ _1104_ VGND VGND 
+ VPWR
+ VPWR _0976_ sky130_fd_sc_hd__a22o_1
X_4581_ net279 _1103_ \cdata[6]\ _1104_ VGND VGND 
+ VPWR
+ VPWR _0975_ sky130_fd_sc_hd__a22o_1
X_4582_ net278 _1103_ \cdata[5]\ _1104_ VGND VGND 
+ VPWR
+ VPWR _0974_ sky130_fd_sc_hd__a22o_1
X_4583_ net277 _1103_ net359 _1104_ VGND VGND 
+ VPWR
+ VPWR _0973_ sky130_fd_sc_hd__a22o_1
X_4584_ net276 _1103_ net361 _1104_ VGND VGND 
+ VPWR
+ VPWR _0972_ sky130_fd_sc_hd__a22o_1
X_4585_ net275 _1103_ net363 _1104_ VGND VGND 
+ VPWR
+ VPWR _0971_ sky130_fd_sc_hd__a22o_1
X_4586_ net299 _1103_ net365 _1104_ VGND VGND 
+ VPWR
+ VPWR _0970_ sky130_fd_sc_hd__a22o_1
X_4587_ net298 _1103_ net367 _1104_ VGND VGND 
+ VPWR
+ VPWR _0969_ sky130_fd_sc_hd__a22o_1
X_4588_ _1040_ _1041_ _0067_ _1030_ VGND VGND 
+ VPWR
+ VPWR _1105_ sky130_fd_sc_hd__or4_4
X_4589_ _1065_ _1105_ VGND VGND VPWR VPWR 
+ _1106_
+ sky130_fd_sc_hd__or2_4
X_4590_ _1023_ _1106_ VGND VGND VPWR VPWR 
+ _1107_
+ sky130_fd_sc_hd__or2_1
X_4591_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__buf_2
X_4592_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__clkinv_2
X_4593_ net297 _1108_ \cdata[7]\ _1109_ VGND VGND 
+ VPWR
+ VPWR _0968_ sky130_fd_sc_hd__a22o_1
X_4594_ net296 _1108_ \cdata[6]\ _1109_ VGND VGND 
+ VPWR
+ VPWR _0967_ sky130_fd_sc_hd__a22o_1
X_4595_ net295 _1108_ \cdata[5]\ _1109_ VGND VGND 
+ VPWR
+ VPWR _0966_ sky130_fd_sc_hd__a22o_1
X_4596_ net294 _1108_ net359 _1109_ VGND VGND 
+ VPWR
+ VPWR _0965_ sky130_fd_sc_hd__a22o_1
X_4597_ net293 _1108_ net361 _1109_ VGND VGND 
+ VPWR
+ VPWR _0964_ sky130_fd_sc_hd__a22o_1
X_4598_ net292 _1108_ net363 _1109_ VGND VGND 
+ VPWR
+ VPWR _0963_ sky130_fd_sc_hd__a22o_1
X_4599_ net285 _1108_ net365 _1109_ VGND VGND 
+ VPWR
+ VPWR _0962_ sky130_fd_sc_hd__a22o_1
X_4600_ net274 _1108_ net367 _1109_ VGND VGND 
+ VPWR
+ VPWR _0961_ sky130_fd_sc_hd__a22o_1
X_4601_ _1028_ _1058_ VGND VGND VPWR VPWR 
+ _1110_
+ sky130_fd_sc_hd__or2_4
X_4602_ _1023_ _1110_ VGND VGND VPWR VPWR 
+ _1111_
+ sky130_fd_sc_hd__or2_1
X_4603_ _1111_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__buf_2
X_4604_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__clkinv_2
X_4605_ net262 _1112_ \cdata[5]\ _1113_ VGND VGND 
+ VPWR
+ VPWR _0960_ sky130_fd_sc_hd__a22o_1
X_4606_ net261 _1112_ net359 _1113_ VGND VGND 
+ VPWR
+ VPWR _0959_ sky130_fd_sc_hd__a22o_1
X_4607_ net260 _1112_ net361 _1113_ VGND VGND 
+ VPWR
+ VPWR _0958_ sky130_fd_sc_hd__a22o_1
X_4608_ net273 _1112_ net363 _1113_ VGND VGND 
+ VPWR
+ VPWR _0957_ sky130_fd_sc_hd__a22o_1
X_4609_ net272 _1112_ net365 _1113_ VGND VGND 
+ VPWR
+ VPWR _0956_ sky130_fd_sc_hd__a22o_1
X_4610_ net271 _1112_ net367 _1113_ VGND VGND 
+ VPWR
+ VPWR _0955_ sky130_fd_sc_hd__a22o_1
X_4611_ _0071_ _0069_ _1029_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1114_ sky130_fd_sc_hd__or4_4
X_4612_ _1028_ _1114_ VGND VGND VPWR VPWR 
+ _1115_
+ sky130_fd_sc_hd__or2_4
X_4613_ _1043_ _1115_ VGND VGND VPWR VPWR 
+ _1116_
+ sky130_fd_sc_hd__or2_1
X_4614_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__clkbuf_2
X_4615_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__inv_2
X_4616_ net269 _1117_ net359 _1118_ VGND VGND 
+ VPWR
+ VPWR _0954_ sky130_fd_sc_hd__a22o_1
X_4617_ net268 _1117_ net361 _1118_ VGND VGND 
+ VPWR
+ VPWR _0953_ sky130_fd_sc_hd__a22o_1
X_4618_ net267 _1117_ net363 _1118_ VGND VGND 
+ VPWR
+ VPWR _0952_ sky130_fd_sc_hd__a22o_1
X_4619_ net266 _1117_ net365 _1118_ VGND VGND 
+ VPWR
+ VPWR _0951_ sky130_fd_sc_hd__a22o_1
X_4620_ net265 _1117_ net367 _1118_ VGND VGND 
+ VPWR
+ VPWR _0950_ sky130_fd_sc_hd__a22o_1
X_4621_ _1040_ _0069_ _0067_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1119_ sky130_fd_sc_hd__or4_4
X_4622_ _1065_ _1119_ VGND VGND VPWR VPWR 
+ _1120_
+ sky130_fd_sc_hd__or2_2
X_4623_ _1043_ _1120_ VGND VGND VPWR VPWR 
+ _1121_
+ sky130_fd_sc_hd__or2_1
X_4624_ net365 net264 _1121_ VGND VGND VPWR 
+ VPWR
+ _1122_ sky130_fd_sc_hd__mux2_1
X_4625_ _1122_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__clkbuf_1
X_4626_ net367 net270 _1121_ VGND VGND VPWR 
+ VPWR
+ _1123_ sky130_fd_sc_hd__mux2_1
X_4627_ _1123_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__clkbuf_1
X_4628_ net375 VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__inv_2
X_4629_ hkspi_disable \gpio_configure[3][3]\ net67 VGND VGND VPWR 
+ VPWR
+ _1125_ sky130_fd_sc_hd__or3_4
X_4630_ _1124_ _1125_ VGND VGND VPWR VPWR 
+ _1126_
+ sky130_fd_sc_hd__nor2_8
X_4631_ _1126_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__buf_12
X_4632_ \hkspi.readmode\ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
X_4633_ \hkspi.state[2]\ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__inv_2
X_4634_ _0154_ _1127_ VGND VGND VPWR VPWR 
+ _1128_
+ sky130_fd_sc_hd__or2_1
X_4635_ _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__clkbuf_4
X_4636_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__inv_2
X_4637_ \hkspi.SDO\ _1129_ _0061_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0947_ sky130_fd_sc_hd__a22o_1
X_4638_ _0261_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__clkbuf_1
X_4639_ _1131_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
X_4640_ \hkspi.ldata[6]\ _1129_ _0060_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0946_ sky130_fd_sc_hd__a22o_1
X_4641_ _0261_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__clkbuf_1
X_4642_ _1132_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
X_4643_ \hkspi.ldata[5]\ _1129_ _0059_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0945_ sky130_fd_sc_hd__a22o_1
X_4644_ _0261_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__clkbuf_1
X_4645_ _1133_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
X_4646_ \hkspi.ldata[4]\ _1129_ _0058_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0944_ sky130_fd_sc_hd__a22o_2
X_4647_ _0261_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__clkbuf_1
X_4648_ _1134_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
X_4649_ \hkspi.ldata[3]\ _1129_ _0057_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0943_ sky130_fd_sc_hd__a22o_1
X_4650_ _0261_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__clkbuf_1
X_4651_ _1135_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
X_4652_ \hkspi.ldata[2]\ _1129_ _0056_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0942_ sky130_fd_sc_hd__a22o_1
X_4653_ _0261_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__clkbuf_1
X_4654_ _1136_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
X_4655_ \hkspi.ldata[1]\ _1129_ _0055_ _1130_ VGND VGND 
+ VPWR
+ VPWR _0941_ sky130_fd_sc_hd__a22o_1
X_4656_ _0261_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__clkbuf_1
X_4657_ _1137_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
X_4658_ \hkspi.count[1]\ \hkspi.count[0]\ \hkspi.count[2]\ VGND VGND VPWR 
+ VPWR
+ _1138_ sky130_fd_sc_hd__or3_2
X_4659_ _1138_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkinv_4
X_4660_ \gpio_configure[17][8]\ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__inv_2
X_4661_ _1036_ _1026_ _1024_ VGND VGND VPWR 
+ VPWR
+ _1140_ sky130_fd_sc_hd__or3_1
X_4662_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__buf_8
X_4663_ _1042_ _1141_ VGND VGND VPWR VPWR 
+ _1142_
+ sky130_fd_sc_hd__or2_4
X_4664_ \gpio_configure[6][0]\ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__clkinv_2
X_4665_ _0073_ _1036_ _1026_ VGND VGND VPWR 
+ VPWR
+ _1144_ sky130_fd_sc_hd__or3_1
X_4666_ _1144_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__buf_8
X_4667_ _1063_ _1145_ VGND VGND VPWR VPWR 
+ _1146_
+ sky130_fd_sc_hd__or2_4
X_4668_ \gpio_configure[7][0]\ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__inv_2
X_4669_ _1040_ _1041_ _0067_ _0065_ VGND VGND 
+ VPWR
+ VPWR _1148_ sky130_fd_sc_hd__or4_4
X_4670_ _1148_ _1145_ VGND VGND VPWR VPWR 
+ _1149_
+ sky130_fd_sc_hd__or2_4
X_4671_ \gpio_configure[35][8]\ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__inv_2
X_4672_ _1031_ _1039_ VGND VGND VPWR VPWR 
+ _1151_
+ sky130_fd_sc_hd__or2_4
X_4673_ _1147_ _1149_ _1150_ _1151_ VGND VGND 
+ VPWR
+ VPWR _1152_ sky130_fd_sc_hd__o22a_1
X_4674_ _1139_ _1142_ _1143_ _1146_ _1152_ VGND 
+ VGND
+ VPWR VPWR _1153_ sky130_fd_sc_hd__o221a_1
X_4675_ \gpio_configure[34][0]\ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__clkinv_2
X_4676_ _1039_ _1114_ VGND VGND VPWR VPWR 
+ _1155_
+ sky130_fd_sc_hd__or2_4
X_4677_ \gpio_configure[2][8]\ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__clkinv_2
X_4678_ _1058_ _1145_ VGND VGND VPWR VPWR 
+ _1157_
+ sky130_fd_sc_hd__or2_4
X_4679_ _1039_ _1089_ VGND VGND VPWR VPWR 
+ _1158_
+ sky130_fd_sc_hd__or2_4
X_4680_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__inv_4
X_4681_ net300 VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__clkinv_4
X_4682_ _1039_ _1100_ VGND VGND VPWR VPWR 
+ _1161_
+ sky130_fd_sc_hd__or2_4
X_4683_ net61 _1159_ _1160_ _1161_ VGND VGND 
+ VPWR
+ VPWR _1162_ sky130_fd_sc_hd__o2bb2a_1
X_4684_ _1154_ _1155_ _1156_ _1157_ _1162_ VGND 
+ VGND
+ VPWR VPWR _1163_ sky130_fd_sc_hd__o221a_1
X_4685_ \gpio_configure[10][8]\ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__inv_2
X_4686_ _1058_ _1141_ VGND VGND VPWR VPWR 
+ _1165_
+ sky130_fd_sc_hd__or2_4
X_4687_ \gpio_configure[4][0]\ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__clkinv_2
X_4688_ _1029_ _0065_ _0071_ _1041_ VGND VGND 
+ VPWR
+ VPWR _1167_ sky130_fd_sc_hd__or4_4
X_4689_ _1167_ _1145_ VGND VGND VPWR VPWR 
+ _1168_
+ sky130_fd_sc_hd__or2_4
X_4690_ \gpio_configure[3][8]\ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__clkinv_4
X_4691_ _1031_ _1145_ VGND VGND VPWR VPWR 
+ _1170_
+ sky130_fd_sc_hd__or2_4
X_4692_ _1169_ _1170_ VGND VGND VPWR VPWR 
+ _1171_
+ sky130_fd_sc_hd__or2_1
X_4693_ _1164_ _1165_ _1166_ _1168_ _1171_ VGND 
+ VGND
+ VPWR VPWR _1172_ sky130_fd_sc_hd__o221a_1
X_4694_ \gpio_configure[8][8]\ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__clkinv_4
X_4695_ _1105_ _1145_ VGND VGND VPWR VPWR 
+ _1174_
+ sky130_fd_sc_hd__or2_4
X_4696_ net36 VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__inv_2
X_4697_ _1039_ _1105_ VGND VGND VPWR VPWR 
+ _1176_
+ sky130_fd_sc_hd__or2_1
X_4698_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__buf_12
X_4699_ \gpio_configure[7][8]\ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__clkinv_2
X_4700_ _1046_ _1145_ VGND VGND VPWR VPWR 
+ _1179_
+ sky130_fd_sc_hd__or2_4
X_4701_ \gpio_configure[5][0]\ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__inv_2
X_4702_ _1119_ _1145_ VGND VGND VPWR VPWR 
+ _1181_
+ sky130_fd_sc_hd__or2_4
X_4703_ _1178_ _1179_ _1180_ _1181_ VGND VGND 
+ VPWR
+ VPWR _1182_ sky130_fd_sc_hd__o22a_1
X_4704_ _1173_ _1174_ _1175_ _1177_ _1182_ VGND 
+ VGND
+ VPWR VPWR _1183_ sky130_fd_sc_hd__o221a_1
X_4705_ _1153_ _1163_ _1172_ _1183_ VGND VGND 
+ VPWR
+ VPWR _1184_ sky130_fd_sc_hd__and4_1
X_4706_ \gpio_configure[14][8]\ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__clkinv_2
X_4707_ _1089_ _1141_ VGND VGND VPWR VPWR 
+ _1186_
+ sky130_fd_sc_hd__or2_4
X_4708_ \gpio_configure[11][0]\ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__inv_2
X_4709_ _1075_ _1141_ VGND VGND VPWR VPWR 
+ _1188_
+ sky130_fd_sc_hd__or2_4
X_4710_ \gpio_configure[15][8]\ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__inv_2
X_4711_ _1046_ _1141_ VGND VGND VPWR VPWR 
+ _1190_
+ sky130_fd_sc_hd__or2_4
X_4712_ \gpio_configure[11][8]\ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__inv_2
X_4713_ _1031_ _1141_ VGND VGND VPWR VPWR 
+ _1192_
+ sky130_fd_sc_hd__or2_4
X_4714_ _1189_ _1190_ _1191_ _1192_ VGND VGND 
+ VPWR
+ VPWR _1193_ sky130_fd_sc_hd__o22a_1
X_4715_ _1185_ _1186_ _1187_ _1188_ _1193_ VGND 
+ VGND
+ VPWR VPWR _1194_ sky130_fd_sc_hd__o221a_1
X_4716_ \gpio_configure[8][0]\ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__clkinv_2
X_4717_ _1100_ _1145_ VGND VGND VPWR VPWR 
+ _1196_
+ sky130_fd_sc_hd__or2_4
X_4718_ \gpio_configure[16][8]\ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__inv_2
X_4719_ _1105_ _1141_ VGND VGND VPWR VPWR 
+ _1198_
+ sky130_fd_sc_hd__or2_4
X_4720_ \gpio_configure[13][0]\ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__clkinv_4
X_4721_ _1119_ _1141_ VGND VGND VPWR VPWR 
+ _1200_
+ sky130_fd_sc_hd__or2_4
X_4722_ \gpio_configure[12][8]\ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__inv_2
X_4723_ _1070_ _1141_ VGND VGND VPWR VPWR 
+ _1202_
+ sky130_fd_sc_hd__or2_4
X_4724_ _1199_ _1200_ _1201_ _1202_ VGND VGND 
+ VPWR
+ VPWR _1203_ sky130_fd_sc_hd__o22a_1
X_4725_ _1195_ _1196_ _1197_ _1198_ _1203_ VGND 
+ VGND
+ VPWR VPWR _1204_ sky130_fd_sc_hd__o221a_1
X_4726_ \gpio_configure[14][0]\ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__clkinv_2
X_4727_ _1063_ _1141_ VGND VGND VPWR VPWR 
+ _1206_
+ sky130_fd_sc_hd__or2_4
X_4728_ \gpio_configure[13][8]\ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__inv_2
X_4729_ _1029_ _1030_ _0071_ _1041_ VGND VGND 
+ VPWR
+ VPWR _1208_ sky130_fd_sc_hd__or4_4
X_4730_ _1208_ _1141_ VGND VGND VPWR VPWR 
+ _1209_
+ sky130_fd_sc_hd__or2_4
X_4731_ _1207_ _1209_ VGND VGND VPWR VPWR 
+ _1210_
+ sky130_fd_sc_hd__or2_1
X_4732_ \gpio_configure[37][0]\ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__inv_2
X_4733_ _1039_ _1119_ VGND VGND VPWR VPWR 
+ _1212_
+ sky130_fd_sc_hd__or2_4
X_4734_ \gpio_configure[10][0]\ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__inv_2
X_4735_ _1114_ _1141_ VGND VGND VPWR VPWR 
+ _1214_
+ sky130_fd_sc_hd__or2_4
X_4736_ _1211_ _1212_ _1213_ _1214_ VGND VGND 
+ VPWR
+ VPWR _1215_ sky130_fd_sc_hd__o22a_1
X_4737_ net71 VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__clkinv_2
X_4738_ _1039_ _1148_ VGND VGND VPWR VPWR 
+ _1217_
+ sky130_fd_sc_hd__or2_1
X_4739_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__buf_6
X_4740_ \gpio_configure[9][0]\ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__clkinv_2
X_4741_ _1053_ _1141_ VGND VGND VPWR VPWR 
+ _1220_
+ sky130_fd_sc_hd__or2_4
X_4742_ \gpio_configure[16][0]\ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__inv_2
X_4743_ _1100_ _1141_ VGND VGND VPWR VPWR 
+ _1222_
+ sky130_fd_sc_hd__or2_4
X_4744_ \gpio_configure[33][0]\ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__inv_2
X_4745_ _1039_ _1053_ VGND VGND VPWR VPWR 
+ _1224_
+ sky130_fd_sc_hd__or2_4
X_4746_ _1221_ _1222_ _1223_ _1224_ VGND VGND 
+ VPWR
+ VPWR _1225_ sky130_fd_sc_hd__o22a_1
X_4747_ _1216_ _1218_ _1219_ _1220_ _1225_ VGND 
+ VGND
+ VPWR VPWR _1226_ sky130_fd_sc_hd__o221a_1
X_4748_ _1205_ _1206_ _1210_ _1215_ _1226_ VGND 
+ VGND
+ VPWR VPWR _1227_ sky130_fd_sc_hd__o2111a_1
X_4749_ \gpio_configure[37][8]\ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__clkinv_2
X_4750_ _1039_ _1208_ VGND VGND VPWR VPWR 
+ _1229_
+ sky130_fd_sc_hd__or2_4
X_4751_ \gpio_configure[35][0]\ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__inv_2
X_4752_ _1039_ _1075_ VGND VGND VPWR VPWR 
+ _1231_
+ sky130_fd_sc_hd__or2_4
X_4753_ hkspi_disable VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__inv_2
X_4754_ net43 VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__inv_2
X_4755_ _1039_ _1046_ VGND VGND VPWR VPWR 
+ _1234_
+ sky130_fd_sc_hd__or2_1
X_4756_ _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__buf_8
X_4757_ _1039_ _1042_ _1232_ _1233_ _1235_ VGND 
+ VGND
+ VPWR VPWR _1236_ sky130_fd_sc_hd__o32a_1
X_4758_ _1228_ _1229_ _1230_ _1231_ _1236_ VGND 
+ VGND
+ VPWR VPWR _1237_ sky130_fd_sc_hd__o221a_1
X_4759_ \gpio_configure[15][0]\ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__clkinv_4
X_4760_ _1148_ _1141_ VGND VGND VPWR VPWR 
+ _1239_
+ sky130_fd_sc_hd__or2_4
X_4761_ \gpio_configure[9][8]\ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__inv_2
X_4762_ _1042_ _1145_ VGND VGND VPWR VPWR 
+ _1241_
+ sky130_fd_sc_hd__or2_4
X_4763_ \gpio_configure[36][8]\ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__inv_2
X_4764_ _1039_ _1070_ VGND VGND VPWR VPWR 
+ _1243_
+ sky130_fd_sc_hd__or2_2
X_4765_ \gpio_configure[4][8]\ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__clkinv_2
X_4766_ _1070_ _1145_ VGND VGND VPWR VPWR 
+ _1245_
+ sky130_fd_sc_hd__or2_4
X_4767_ _1242_ _1243_ _1244_ _1245_ VGND VGND 
+ VPWR
+ VPWR _1246_ sky130_fd_sc_hd__o22a_1
X_4768_ _1238_ _1239_ _1240_ _1241_ _1246_ VGND 
+ VGND
+ VPWR VPWR _1247_ sky130_fd_sc_hd__o221a_1
X_4769_ \gpio_configure[1][0]\ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__inv_2
X_4770_ _1053_ _1145_ VGND VGND VPWR VPWR 
+ _1249_
+ sky130_fd_sc_hd__or2_4
X_4771_ \gpio_configure[36][0]\ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__inv_2
X_4772_ _1039_ _1167_ VGND VGND VPWR VPWR 
+ _1251_
+ sky130_fd_sc_hd__or2_4
X_4773_ \gpio_configure[2][0]\ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__inv_2
X_4774_ _1114_ _1145_ VGND VGND VPWR VPWR 
+ _1253_
+ sky130_fd_sc_hd__or2_4
X_4775_ \gpio_configure[6][8]\ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__clkinv_2
X_4776_ _1089_ _1145_ VGND VGND VPWR VPWR 
+ _1255_
+ sky130_fd_sc_hd__or2_4
X_4777_ _1252_ _1253_ _1254_ _1255_ VGND VGND 
+ VPWR
+ VPWR _1256_ sky130_fd_sc_hd__o22a_2
X_4778_ _1248_ _1249_ _1250_ _1251_ _1256_ VGND 
+ VGND
+ VPWR VPWR _1257_ sky130_fd_sc_hd__o221a_1
X_4779_ \gpio_configure[12][0]\ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__clkinv_2
X_4780_ _1167_ _1141_ VGND VGND VPWR VPWR 
+ _1259_
+ sky130_fd_sc_hd__or2_4
X_4781_ net52 VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__clkinv_2
X_4782_ _1039_ _1063_ VGND VGND VPWR VPWR 
+ _1261_
+ sky130_fd_sc_hd__or2_1
X_4783_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__buf_12
X_4784_ \gpio_configure[5][8]\ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__inv_2
X_4785_ _1208_ _1145_ VGND VGND VPWR VPWR 
+ _1264_
+ sky130_fd_sc_hd__or2_4
X_4786_ \gpio_configure[34][8]\ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__inv_2
X_4787_ _1039_ _1058_ VGND VGND VPWR VPWR 
+ _1266_
+ sky130_fd_sc_hd__or2_4
X_4788_ _1263_ _1264_ _1265_ _1266_ VGND VGND 
+ VPWR
+ VPWR _1267_ sky130_fd_sc_hd__o22a_2
X_4789_ _1258_ _1259_ _1260_ _1262_ _1267_ VGND 
+ VGND
+ VPWR VPWR _1268_ sky130_fd_sc_hd__o221a_1
X_4790_ _1237_ _1247_ _1257_ _1268_ VGND VGND 
+ VPWR
+ VPWR _1269_ sky130_fd_sc_hd__and4_1
X_4791_ _1194_ _1204_ _1227_ _1269_ VGND VGND 
+ VPWR
+ VPWR _1270_ sky130_fd_sc_hd__and4_1
X_4792_ net281 VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__inv_2
X_4793_ \gpio_configure[27][0]\ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__clkinv_4
X_4794_ _1052_ _1075_ VGND VGND VPWR VPWR 
+ _1273_
+ sky130_fd_sc_hd__or2_4
X_4795_ \gpio_configure[0][8]\ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__inv_2
X_4796_ _1028_ _1105_ VGND VGND VPWR VPWR 
+ _1275_
+ sky130_fd_sc_hd__or2_4
X_4797_ net265 VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__inv_2
X_4798_ _1274_ _1275_ _1276_ _1115_ VGND VGND 
+ VPWR
+ VPWR _1277_ sky130_fd_sc_hd__o22a_1
X_4799_ _1271_ _1096_ _1272_ _1273_ _1277_ VGND 
+ VGND
+ VPWR VPWR _1278_ sky130_fd_sc_hd__o221a_1
X_4800_ \gpio_configure[24][8]\ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__clkinv_2
X_4801_ _0073_ _0075_ _1037_ VGND VGND VPWR 
+ VPWR
+ _1280_ sky130_fd_sc_hd__or3_1
X_4802_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__buf_6
X_4803_ _1105_ _1281_ VGND VGND VPWR VPWR 
+ _1282_
+ sky130_fd_sc_hd__or2_4
X_4804_ \gpio_configure[17][0]\ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__clkinv_4
X_4805_ _1053_ _1281_ VGND VGND VPWR VPWR 
+ _1284_
+ sky130_fd_sc_hd__or2_4
X_4806_ reset_reg \hkspi.pre_pass_thru_mgmt\ \hkspi.pass_thru_mgmt_delay\ VGND VGND VPWR 
+ VPWR
+ _1285_ sky130_fd_sc_hd__or3_1
X_4807_ _1285_ VGND VGND VPWR VPWR net304 sky130_fd_sc_hd__buf_2
X_4808_ net304 VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__inv_2
X_4809_ \gpio_configure[25][8]\ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__clkinv_2
X_4810_ _1042_ _1281_ VGND VGND VPWR VPWR 
+ _1288_
+ sky130_fd_sc_hd__or2_4
X_4811_ _1046_ _1065_ _1286_ _1287_ _1288_ VGND 
+ VGND
+ VPWR VPWR _1289_ sky130_fd_sc_hd__o32a_1
X_4812_ _1279_ _1282_ _1283_ _1284_ _1289_ VGND 
+ VGND
+ VPWR VPWR _1290_ sky130_fd_sc_hd__o221a_1
X_4813_ net325 VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__inv_2
X_4814_ \gpio_configure[26][0]\ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__inv_6
X_4815_ _1052_ _1114_ VGND VGND VPWR VPWR 
+ _1293_
+ sky130_fd_sc_hd__or2_4
X_4816_ \gpio_configure[31][0]\ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__inv_4
X_4817_ _1052_ _1148_ VGND VGND VPWR VPWR 
+ _1295_
+ sky130_fd_sc_hd__or2_4
X_4818_ net270 VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__clkinv_2
X_4819_ _1294_ _1295_ _1296_ _1120_ VGND VGND 
+ VPWR
+ VPWR _1297_ sky130_fd_sc_hd__o22a_1
X_4820_ _1291_ _1076_ _1292_ _1293_ _1297_ VGND 
+ VGND
+ VPWR VPWR _1298_ sky130_fd_sc_hd__o221a_1
X_4821_ net20 VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__inv_2
X_4822_ _1065_ _1075_ VGND VGND VPWR VPWR 
+ _1300_
+ sky130_fd_sc_hd__or2_4
X_4823_ \gpio_configure[1][8]\ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__inv_2
X_4824_ _1028_ _1042_ VGND VGND VPWR VPWR 
+ _1302_
+ sky130_fd_sc_hd__or2_4
X_4825_ irq_1_inputsrc VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__inv_2
X_4826_ _1028_ _1148_ VGND VGND VPWR VPWR 
+ _1304_
+ sky130_fd_sc_hd__or2_1
X_4827_ serial_busy VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__clkinv_2
X_4828_ _1303_ _1304_ _1305_ _1032_ VGND VGND 
+ VPWR
+ VPWR _1306_ sky130_fd_sc_hd__o22a_1
X_4829_ _1299_ _1300_ _1301_ _1302_ _1306_ VGND 
+ VGND
+ VPWR VPWR _1307_ sky130_fd_sc_hd__o221a_1
X_4830_ _1278_ _1290_ _1298_ _1307_ VGND VGND 
+ VPWR
+ VPWR _1308_ sky130_fd_sc_hd__and4_1
X_4831_ net109 VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__clkinv_2
X_4832_ _1028_ _1167_ VGND VGND VPWR VPWR 
+ _1310_
+ sky130_fd_sc_hd__or2_4
X_4833_ \gpio_configure[32][0]\ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__inv_4
X_4834_ _1052_ _1100_ VGND VGND VPWR VPWR 
+ _1312_
+ sky130_fd_sc_hd__or2_4
X_4835_ trap_output_dest VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__clkinv_4
X_4836_ \gpio_configure[27][8]\ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__clkinv_2
X_4837_ _1031_ _1052_ VGND VGND VPWR VPWR 
+ _1315_
+ sky130_fd_sc_hd__or2_4
X_4838_ _1313_ _1047_ _1314_ _1315_ VGND VGND 
+ VPWR
+ VPWR _1316_ sky130_fd_sc_hd__o22a_1
X_4839_ _1309_ _1310_ _1311_ _1312_ _1316_ VGND 
+ VGND
+ VPWR VPWR _1317_ sky130_fd_sc_hd__o221a_1
X_4840_ net100 VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__clkinv_2
X_4841_ _1028_ _1208_ VGND VGND VPWR VPWR 
+ _1319_
+ sky130_fd_sc_hd__or2_4
X_4842_ \gpio_configure[3][0]\ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__clkinv_4
X_4843_ _1075_ _1145_ VGND VGND VPWR VPWR 
+ _1321_
+ sky130_fd_sc_hd__or2_4
X_4844_ _1031_ _1065_ VGND VGND VPWR VPWR 
+ _1322_
+ sky130_fd_sc_hd__or2_1
X_4845_ _1318_ _1319_ _1320_ _1321_ _1322_ VGND 
+ VGND
+ VPWR VPWR _1323_ sky130_fd_sc_hd__o221a_1
X_4846_ \gpio_configure[24][0]\ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__inv_2
X_4847_ _1100_ _1281_ VGND VGND VPWR VPWR 
+ _1325_
+ sky130_fd_sc_hd__or2_4
X_4848_ \gpio_configure[20][8]\ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__clkinv_2
X_4849_ _1070_ _1281_ VGND VGND VPWR VPWR 
+ _1327_
+ sky130_fd_sc_hd__or2_4
X_4850_ \gpio_configure[30][0]\ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__inv_2
X_4851_ _1052_ _1063_ VGND VGND VPWR VPWR 
+ _1329_
+ sky130_fd_sc_hd__or2_4
X_4852_ net316 VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__inv_2
X_4853_ _1328_ _1329_ _1330_ _1071_ VGND VGND 
+ VPWR
+ VPWR _1331_ sky130_fd_sc_hd__o22a_1
X_4854_ _1324_ _1325_ _1326_ _1327_ _1331_ VGND 
+ VGND
+ VPWR VPWR _1332_ sky130_fd_sc_hd__o221a_1
X_4855_ \gpio_configure[29][0]\ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__inv_2
X_4856_ _1052_ _1119_ VGND VGND VPWR VPWR 
+ _1334_
+ sky130_fd_sc_hd__or2_4
X_4857_ \gpio_configure[25][0]\ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__inv_2
X_4858_ \gpio_configure[31][8]\ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__inv_2
X_4859_ _1046_ _1052_ VGND VGND VPWR VPWR 
+ _1337_
+ sky130_fd_sc_hd__or2_4
X_4860_ net93 VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__inv_2
X_4861_ _1028_ _1089_ VGND VGND VPWR VPWR 
+ _1339_
+ sky130_fd_sc_hd__or2_4
X_4862_ _1336_ _1337_ _1338_ _1339_ VGND VGND 
+ VPWR
+ VPWR _1340_ sky130_fd_sc_hd__o22a_1
X_4863_ _1333_ _1334_ _1335_ _1054_ _1340_ VGND 
+ VGND
+ VPWR VPWR _1341_ sky130_fd_sc_hd__o221a_1
X_4864_ _1317_ _1323_ _1332_ _1341_ VGND VGND 
+ VPWR
+ VPWR _1342_ sky130_fd_sc_hd__and4_1
X_4865_ \gpio_configure[30][8]\ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__clkinv_4
X_4866_ _1052_ _1089_ VGND VGND VPWR VPWR 
+ _1344_
+ sky130_fd_sc_hd__or2_4
X_4867_ net130 VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__inv_4
X_4868_ _1028_ _1063_ VGND VGND VPWR VPWR 
+ _1346_
+ sky130_fd_sc_hd__or2_4
X_4869_ net4 VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__inv_2
X_4870_ _1065_ _1208_ VGND VGND VPWR VPWR 
+ _1348_
+ sky130_fd_sc_hd__or2_4
X_4871_ net290 VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__inv_2
X_4872_ _1347_ _1348_ _1349_ _1092_ VGND VGND 
+ VPWR
+ VPWR _1350_ sky130_fd_sc_hd__o22a_2
X_4873_ _1343_ _1344_ _1345_ _1346_ _1350_ VGND 
+ VGND
+ VPWR VPWR _1351_ sky130_fd_sc_hd__o221a_1
X_4874_ net271 VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__inv_2
X_4875_ \gpio_configure[0][0]\ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__inv_2
X_4876_ _1028_ _1100_ VGND VGND VPWR VPWR 
+ _1353_
+ sky130_fd_sc_hd__or2_4
X_4877_ \gpio_configure[18][0]\ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__inv_2
X_4878_ _1114_ _1281_ VGND VGND VPWR VPWR 
+ _1355_
+ sky130_fd_sc_hd__or2_4
X_4879_ net204 VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__inv_2
X_4880_ _1354_ _1355_ _1356_ _1066_ VGND VGND 
+ VPWR
+ VPWR _1357_ sky130_fd_sc_hd__o22a_2
X_4881_ _1352_ _1110_ _0099_ _1353_ _1357_ VGND 
+ VGND
+ VPWR VPWR _1358_ sky130_fd_sc_hd__o221a_1
X_4882_ \gpio_configure[26][8]\ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__inv_2
X_4883_ \gpio_configure[28][8]\ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__inv_2
X_4884_ _1052_ _1070_ VGND VGND VPWR VPWR 
+ _1361_
+ sky130_fd_sc_hd__or2_4
X_4885_ _1065_ _1167_ net34 VGND VGND VPWR 
+ VPWR
+ _1362_ sky130_fd_sc_hd__or3b_1
X_4886_ _1359_ _1059_ _1360_ _1361_ _1362_ VGND 
+ VGND
+ VPWR VPWR _1363_ sky130_fd_sc_hd__o221a_1
X_4887_ net274 VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__inv_2
X_4888_ \gpio_configure[29][8]\ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__inv_2
X_4889_ _1052_ _1208_ VGND VGND VPWR VPWR 
+ _1366_
+ sky130_fd_sc_hd__or2_4
X_4890_ \gpio_configure[33][8]\ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__inv_2
X_4891_ _1042_ _1052_ VGND VGND VPWR VPWR 
+ _1368_
+ sky130_fd_sc_hd__or2_4
X_4892_ net123 VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__inv_2
X_4893_ _1028_ _1119_ VGND VGND VPWR VPWR 
+ _1370_
+ sky130_fd_sc_hd__or2_4
X_4894_ _1367_ _1368_ _1369_ _1370_ VGND VGND 
+ VPWR
+ VPWR _1371_ sky130_fd_sc_hd__o22a_1
X_4895_ _1364_ _1106_ _1365_ _1366_ _1371_ VGND 
+ VGND
+ VPWR VPWR _1372_ sky130_fd_sc_hd__o221a_1
X_4896_ _1351_ _1358_ _1363_ _1372_ VGND VGND 
+ VPWR
+ VPWR _1373_ sky130_fd_sc_hd__and4_1
X_4897_ \gpio_configure[22][0]\ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__clkinv_4
X_4898_ _1063_ _1281_ VGND VGND VPWR VPWR 
+ _1375_
+ sky130_fd_sc_hd__or2_4
X_4899_ \gpio_configure[21][8]\ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__clkinv_2
X_4900_ _1281_ _1208_ VGND VGND VPWR VPWR 
+ _1377_
+ sky130_fd_sc_hd__or2_4
X_4901_ net125 VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__inv_2
X_4902_ \gpio_configure[32][8]\ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__inv_2
X_4903_ _1052_ _1105_ VGND VGND VPWR VPWR 
+ _1380_
+ sky130_fd_sc_hd__or2_4
X_4904_ _1065_ _1148_ _1378_ _1379_ _1380_ VGND 
+ VGND
+ VPWR VPWR _1381_ sky130_fd_sc_hd__o32a_1
X_4905_ _1374_ _1375_ _1376_ _1377_ _1381_ VGND 
+ VGND
+ VPWR VPWR _1382_ sky130_fd_sc_hd__o221a_1
X_4906_ net11 VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__inv_2
X_4907_ _1065_ _1070_ VGND VGND VPWR VPWR 
+ _1384_
+ sky130_fd_sc_hd__or2_4
X_4908_ net298 VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__inv_2
X_4909_ net263 VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__inv_2
X_4910_ \gpio_configure[28][0]\ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__inv_4
X_4911_ _1052_ _1167_ VGND VGND VPWR VPWR 
+ _1388_
+ sky130_fd_sc_hd__or2_4
X_4912_ _1065_ _1089_ _1386_ _1387_ _1388_ VGND 
+ VGND
+ VPWR VPWR _1389_ sky130_fd_sc_hd__o32a_1
X_4913_ _1383_ _1384_ _1385_ _1101_ _1389_ VGND 
+ VGND
+ VPWR VPWR _1390_ sky130_fd_sc_hd__o221a_2
X_4914_ \gpio_configure[20][0]\ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__clkinv_2
X_4915_ _1167_ _1281_ VGND VGND VPWR VPWR 
+ _1392_
+ sky130_fd_sc_hd__or2_4
X_4916_ \gpio_configure[21][0]\ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__inv_2
X_4917_ _1119_ _1281_ VGND VGND VPWR VPWR 
+ _1394_
+ sky130_fd_sc_hd__or2_4
X_4918_ \gpio_configure[19][8]\ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__clkinv_2
X_4919_ _1031_ _1281_ VGND VGND VPWR VPWR 
+ _1396_
+ sky130_fd_sc_hd__or2_4
X_4920_ \gpio_configure[18][8]\ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__clkinv_2
X_4921_ _1058_ _1281_ VGND VGND VPWR VPWR 
+ _1398_
+ sky130_fd_sc_hd__or2_4
X_4922_ _1395_ _1396_ _1397_ _1398_ VGND VGND 
+ VPWR
+ VPWR _1399_ sky130_fd_sc_hd__o22a_2
X_4923_ _1391_ _1392_ _1393_ _1394_ _1399_ VGND 
+ VGND
+ VPWR VPWR _1400_ sky130_fd_sc_hd__o221a_1
X_4924_ \gpio_configure[22][8]\ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__clkinv_2
X_4925_ _1089_ _1281_ VGND VGND VPWR VPWR 
+ _1402_
+ sky130_fd_sc_hd__or2_4
X_4926_ \gpio_configure[23][0]\ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__clkinv_4
X_4927_ _1148_ _1281_ VGND VGND VPWR VPWR 
+ _1404_
+ sky130_fd_sc_hd__or2_4
X_4928_ \gpio_configure[19][0]\ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__inv_2
X_4929_ _1075_ _1281_ VGND VGND VPWR VPWR 
+ _1406_
+ sky130_fd_sc_hd__or2_4
X_4930_ \gpio_configure[23][8]\ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__clkinv_2
X_4931_ _1046_ _1281_ VGND VGND VPWR VPWR 
+ _1408_
+ sky130_fd_sc_hd__or2_4
X_4932_ _1405_ _1406_ _1407_ _1408_ VGND VGND 
+ VPWR
+ VPWR _1409_ sky130_fd_sc_hd__o22a_1
X_4933_ _1401_ _1402_ _1403_ _1404_ _1409_ VGND 
+ VGND
+ VPWR VPWR _1410_ sky130_fd_sc_hd__o221a_1
X_4934_ _1382_ _1390_ _1400_ _1410_ VGND VGND 
+ VPWR
+ VPWR _1411_ sky130_fd_sc_hd__and4_1
X_4935_ _1308_ _1342_ _1373_ _1411_ VGND VGND 
+ VPWR
+ VPWR _1412_ sky130_fd_sc_hd__and4_2
X_4936_ _1184_ _1270_ _1412_ VGND VGND VPWR 
+ VPWR
+ _1413_ sky130_fd_sc_hd__nand3_4
X_4937_ _1130_ _0062_ _1413_ \hkspi.ldata[0]\ _1129_ VGND 
+ VGND
+ VPWR VPWR _0940_ sky130_fd_sc_hd__a32o_1
X_4938_ _0261_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__clkbuf_1
X_4939_ _1414_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
X_4940_ \hkspi.count[2]\ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__inv_2
X_4941_ \hkspi.count[1]\ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__inv_2
X_4942_ \hkspi.count[0]\ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__clkinv_2
X_4943_ _1415_ _1416_ _1417_ VGND VGND VPWR 
+ VPWR
+ _1418_ sky130_fd_sc_hd__or3_1
X_4944_ _1418_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__clkbuf_4
X_4945_ _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__clkinv_2
X_4946_ \hkspi.wrstb\ \hkspi.writemode\ \hkspi.state[2]\ _1420_ VGND VGND 
+ VPWR
+ VPWR _0939_ sky130_fd_sc_hd__o211a_1
X_4947_ _0261_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__clkbuf_1
X_4948_ _1421_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
X_4949_ net58 VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__clkinv_2
X_4950_ \hkspi.count[2]\ \hkspi.count[1]\ _1417_ VGND VGND VPWR 
+ VPWR
+ _1423_ sky130_fd_sc_hd__and3_1
X_4951_ \hkspi.state[0]\ _1423_ VGND VGND VPWR VPWR 
+ _1424_
+ sky130_fd_sc_hd__nand2_1
X_4952_ \hkspi.pre_pass_thru_user\ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__inv_2
X_4953_ \hkspi.pre_pass_thru_mgmt\ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__inv_2
X_4954_ _1426_ _1419_ \hkspi.count[2]\ \hkspi.state[0]\ \hkspi.count[1]\ VGND 
+ VGND
+ VPWR VPWR _1427_ sky130_fd_sc_hd__o2111a_1
X_4955_ _1422_ _1424_ _1425_ _1427_ VGND VGND 
+ VPWR
+ VPWR _0938_ sky130_fd_sc_hd__o22ai_1
X_4956_ _0261_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__clkbuf_1
X_4957_ _1428_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
X_4958_ \hkspi.count[1]\ _1417_ VGND VGND VPWR VPWR 
+ _1429_
+ sky130_fd_sc_hd__nor2_1
X_4959_ \hkspi.state[0]\ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkinv_4
X_4960_ _1415_ _0087_ _1417_ \hkspi.pre_pass_thru_mgmt\ VGND VGND 
+ VPWR
+ VPWR _1430_ sky130_fd_sc_hd__o31a_1
X_4961_ \hkspi.count[2]\ \hkspi.state[0]\ net58 _1429_ _1430_ VGND 
+ VGND
+ VPWR VPWR _0937_ sky130_fd_sc_hd__a41o_1
X_4962_ _0261_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__clkbuf_1
X_4963_ _1431_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
X_4964_ \hkspi.state[0]\ _1127_ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _1432_ sky130_fd_sc_hd__or3_1
X_4965_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__buf_8
X_4966_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__clkinv_2
X_4967_ \hkspi.odata[7]\ _1433_ \hkspi.odata[6]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0936_ sky130_fd_sc_hd__a22o_1
X_4968_ _0261_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__clkbuf_1
X_4969_ _1435_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
X_4970_ \hkspi.odata[6]\ _1433_ \hkspi.odata[5]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0935_ sky130_fd_sc_hd__a22o_1
X_4971_ _0261_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__clkbuf_1
X_4972_ _1436_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
X_4973_ \hkspi.odata[5]\ _1433_ \hkspi.odata[4]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0934_ sky130_fd_sc_hd__a22o_1
X_4974_ _0261_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__clkbuf_1
X_4975_ _1437_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
X_4976_ \hkspi.odata[4]\ _1433_ \hkspi.odata[3]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0933_ sky130_fd_sc_hd__a22o_1
X_4977_ _0261_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__clkbuf_1
X_4978_ _1438_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
X_4979_ \hkspi.odata[3]\ _1433_ \hkspi.odata[2]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0932_ sky130_fd_sc_hd__a22o_1
X_4980_ _0261_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__clkbuf_1
X_4981_ _1439_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
X_4982_ \hkspi.odata[2]\ _1433_ \hkspi.odata[1]\ _1434_ VGND VGND 
+ VPWR
+ VPWR _0931_ sky130_fd_sc_hd__a22o_1
X_4983_ _0261_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__clkbuf_1
X_4984_ _1440_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
X_4985_ \hkspi.odata[1]\ _1433_ net58 _1434_ VGND VGND 
+ VPWR
+ VPWR _0930_ sky130_fd_sc_hd__a22o_1
X_4986_ _0261_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__clkbuf_1
X_4987_ _1441_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
X_4988_ \hkspi.fixed[2]\ \hkspi.fixed[1]\ VGND VGND VPWR VPWR 
+ _1442_
+ sky130_fd_sc_hd__nor2_1
X_4989_ \hkspi.count[1]\ \hkspi.count[0]\ \hkspi.count[2]\ VGND VGND VPWR 
+ VPWR
+ _1443_ sky130_fd_sc_hd__o21a_1
X_4990_ _1419_ _1442_ _1433_ _0087_ _1443_ VGND 
+ VGND
+ VPWR VPWR _1444_ sky130_fd_sc_hd__o32a_1
X_4991_ _1444_ _0090_ VGND VGND VPWR VPWR 
+ _1445_
+ sky130_fd_sc_hd__or2b_1
X_4992_ _0045_ \hkspi.fixed[2]\ _1445_ VGND VGND VPWR 
+ VPWR
+ _1446_ sky130_fd_sc_hd__mux2_1
X_4993_ _1446_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__clkbuf_1
X_4994_ _0261_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__clkbuf_1
X_4995_ _1447_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
X_4996_ _0044_ \hkspi.fixed[1]\ _1445_ VGND VGND VPWR 
+ VPWR
+ _1448_ sky130_fd_sc_hd__mux2_1
X_4997_ _1448_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__clkbuf_1
X_4998_ _1126_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__buf_8
X_4999_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__clkbuf_1
X_5000_ _1450_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
X_5001_ _0043_ \hkspi.fixed[0]\ _1445_ VGND VGND VPWR 
+ VPWR
+ _1451_ sky130_fd_sc_hd__mux2_1
X_5002_ _1451_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_1
X_5003_ _1449_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__clkbuf_1
X_5004_ _1452_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
X_5005_ \hkspi.count[1]\ _1417_ \hkspi.count[2]\ _0087_ VGND VGND 
+ VPWR
+ VPWR _1453_ sky130_fd_sc_hd__or4_1
X_5006_ _1453_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_5007_ net58 \hkspi.readmode\ _0089_ VGND VGND VPWR 
+ VPWR
+ _1454_ sky130_fd_sc_hd__mux2_1
X_5008_ _1454_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__clkbuf_1
X_5009_ _1449_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__clkbuf_1
X_5010_ _1455_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
X_5011_ _0087_ _1138_ VGND VGND VPWR VPWR 
+ _1456_
+ sky130_fd_sc_hd__or2_1
X_5012_ \hkspi.state[0]\ _0062_ net58 \hkspi.writemode\ _1456_ VGND 
+ VGND
+ VPWR VPWR _0925_ sky130_fd_sc_hd__a32o_1
X_5013_ _1023_ _1181_ VGND VGND VPWR VPWR 
+ _1457_
+ sky130_fd_sc_hd__or2_1
X_5014_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__buf_2
X_5015_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__inv_2
X_5016_ \gpio_configure[5][7]\ _1458_ \cdata[7]\ _1459_ VGND VGND 
+ VPWR
+ VPWR _0924_ sky130_fd_sc_hd__a22o_1
X_5017_ \gpio_configure[5][6]\ _1458_ \cdata[6]\ _1459_ VGND VGND 
+ VPWR
+ VPWR _0923_ sky130_fd_sc_hd__a22o_1
X_5018_ \gpio_configure[5][5]\ _1458_ \cdata[5]\ _1459_ VGND VGND 
+ VPWR
+ VPWR _0922_ sky130_fd_sc_hd__a22o_1
X_5019_ \gpio_configure[5][4]\ _1458_ net360 _1459_ VGND VGND 
+ VPWR
+ VPWR _0921_ sky130_fd_sc_hd__a22o_1
X_5020_ \gpio_configure[5][3]\ _1458_ net362 _1459_ VGND VGND 
+ VPWR
+ VPWR _0920_ sky130_fd_sc_hd__a22o_1
X_5021_ \gpio_configure[5][2]\ _1458_ net364 _1459_ VGND VGND 
+ VPWR
+ VPWR _0919_ sky130_fd_sc_hd__a22o_1
X_5022_ \gpio_configure[5][1]\ _1458_ net366 _1459_ VGND VGND 
+ VPWR
+ VPWR _0918_ sky130_fd_sc_hd__a22o_1
X_5023_ \gpio_configure[5][0]\ _1458_ net368 _1459_ VGND VGND 
+ VPWR
+ VPWR _0917_ sky130_fd_sc_hd__a22o_1
X_5024_ _1043_ _1170_ VGND VGND VPWR VPWR 
+ _1460_
+ sky130_fd_sc_hd__or2_2
X_5025_ _1460_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__clkbuf_2
X_5026_ _1461_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__inv_2
X_5027_ \gpio_configure[3][12]\ _1461_ net360 _1462_ VGND VGND 
+ VPWR
+ VPWR _0916_ sky130_fd_sc_hd__a22o_1
X_5028_ \gpio_configure[3][11]\ _1461_ \cdata[3]\ _1462_ VGND VGND 
+ VPWR
+ VPWR _0915_ sky130_fd_sc_hd__a22o_1
X_5029_ \gpio_configure[3][10]\ _1461_ \cdata[2]\ _1462_ VGND VGND 
+ VPWR
+ VPWR _0914_ sky130_fd_sc_hd__a22o_1
X_5030_ \gpio_configure[3][9]\ _1461_ \cdata[1]\ _1462_ VGND VGND 
+ VPWR
+ VPWR _0913_ sky130_fd_sc_hd__a22o_1
X_5031_ \gpio_configure[3][8]\ _1461_ \cdata[0]\ _1462_ VGND VGND 
+ VPWR
+ VPWR _0912_ sky130_fd_sc_hd__a22o_1
X_5032_ _1449_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__clkbuf_1
X_5033_ _1463_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
X_5034_ \hkspi.state[4]\ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__inv_2
X_5035_ \hkspi.state[0]\ \hkspi.state[2]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _1465_ sky130_fd_sc_hd__or3_1
X_5036_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__inv_2
X_5037_ \hkspi.state[1]\ _1464_ _1466_ \hkspi.pass_thru_user\ VGND VGND 
+ VPWR
+ VPWR _0911_ sky130_fd_sc_hd__a31o_1
X_5038_ _4407_ _1086_ \wbbd_addr[6]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0910_ sky130_fd_sc_hd__a22o_1
X_5039_ _4406_ _1086_ \wbbd_addr[5]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0909_ sky130_fd_sc_hd__a22o_1
X_5040_ _4405_ _1086_ \wbbd_addr[4]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0908_ sky130_fd_sc_hd__a22o_1
X_5041_ _4404_ _1086_ \wbbd_addr[3]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0907_ sky130_fd_sc_hd__a22o_1
X_5042_ _4403_ _1086_ \wbbd_addr[2]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0906_ sky130_fd_sc_hd__a22o_1
X_5043_ _4402_ _1086_ \wbbd_addr[1]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0905_ sky130_fd_sc_hd__a22o_1
X_5044_ _4401_ _1086_ \wbbd_addr[0]\ _1087_ VGND VGND 
+ VPWR
+ VPWR _0904_ sky130_fd_sc_hd__a22o_1
X_5045_ _1023_ _1253_ VGND VGND VPWR VPWR 
+ _1467_
+ sky130_fd_sc_hd__or2_1
X_5046_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__clkbuf_4
X_5047_ _1468_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__inv_2
X_5048_ \gpio_configure[2][7]\ _1468_ \cdata[7]\ _1469_ VGND VGND 
+ VPWR
+ VPWR _0903_ sky130_fd_sc_hd__a22o_1
X_5049_ \gpio_configure[2][6]\ _1468_ \cdata[6]\ _1469_ VGND VGND 
+ VPWR
+ VPWR _0902_ sky130_fd_sc_hd__a22o_1
X_5050_ \gpio_configure[2][5]\ _1468_ \cdata[5]\ _1469_ VGND VGND 
+ VPWR
+ VPWR _0901_ sky130_fd_sc_hd__a22o_1
X_5051_ \gpio_configure[2][4]\ _1468_ net360 _1469_ VGND VGND 
+ VPWR
+ VPWR _0900_ sky130_fd_sc_hd__a22o_1
X_5052_ \gpio_configure[2][3]\ _1468_ net362 _1469_ VGND VGND 
+ VPWR
+ VPWR _0899_ sky130_fd_sc_hd__a22o_1
X_5053_ \gpio_configure[2][2]\ _1468_ net364 _1469_ VGND VGND 
+ VPWR
+ VPWR _0898_ sky130_fd_sc_hd__a22o_1
X_5054_ \gpio_configure[2][1]\ _1468_ net366 _1469_ VGND VGND 
+ VPWR
+ VPWR _0897_ sky130_fd_sc_hd__a22o_1
X_5055_ \gpio_configure[2][0]\ _1468_ net368 _1469_ VGND VGND 
+ VPWR
+ VPWR _0896_ sky130_fd_sc_hd__a22o_1
X_5056_ net199 net202 _1082_ VGND VGND VPWR 
+ VPWR
+ _1470_ sky130_fd_sc_hd__a21oi_1
X_5057_ net202 net200 _1084_ VGND VGND VPWR 
+ VPWR
+ _1471_ sky130_fd_sc_hd__a21oi_1
X_5058_ net202 net198 VGND VGND VPWR VPWR 
+ _1472_
+ sky130_fd_sc_hd__and2_1
X_5059_ net202 net197 VGND VGND VPWR VPWR 
+ _1473_
+ sky130_fd_sc_hd__and2_1
X_5060_ _1473_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
X_5061_ _1083_ _1472_ _1081_ _0088_ VGND VGND 
+ VPWR
+ VPWR _1474_ sky130_fd_sc_hd__o22ai_1
X_5062_ _1470_ _1471_ _1474_ _1087_ VGND VGND 
+ VPWR
+ VPWR _1475_ sky130_fd_sc_hd__or4_1
X_5063_ _1475_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__clkbuf_4
X_5064_ _4400_ \wbbd_data[7]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1477_ sky130_fd_sc_hd__mux2_1
X_5065_ _1477_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__clkbuf_1
X_5066_ _4399_ \wbbd_data[6]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1478_ sky130_fd_sc_hd__mux2_1
X_5067_ _1478_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__clkbuf_1
X_5068_ _4398_ \wbbd_data[5]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1479_ sky130_fd_sc_hd__mux2_1
X_5069_ _1479_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__clkbuf_1
X_5070_ _4397_ \wbbd_data[4]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1480_ sky130_fd_sc_hd__mux2_1
X_5071_ _1480_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__clkbuf_1
X_5072_ _4396_ \wbbd_data[3]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1481_ sky130_fd_sc_hd__mux2_1
X_5073_ _1481_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__clkbuf_1
X_5074_ _4395_ \wbbd_data[2]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1482_ sky130_fd_sc_hd__mux2_1
X_5075_ _1482_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__clkbuf_1
X_5076_ _4394_ \wbbd_data[1]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1483_ sky130_fd_sc_hd__mux2_1
X_5077_ _1483_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__clkbuf_1
X_5078_ _4393_ \wbbd_data[0]\ _1476_ VGND VGND VPWR 
+ VPWR
+ _1484_ sky130_fd_sc_hd__mux2_1
X_5079_ _1484_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__clkbuf_1
X_5080_ _1043_ _1157_ VGND VGND VPWR VPWR 
+ _1485_
+ sky130_fd_sc_hd__or2_1
X_5081_ _1485_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__clkbuf_2
X_5082_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__inv_2
X_5083_ \gpio_configure[2][12]\ _1486_ net359 _1487_ VGND VGND 
+ VPWR
+ VPWR _0887_ sky130_fd_sc_hd__a22o_1
X_5084_ \gpio_configure[2][11]\ _1486_ net361 _1487_ VGND VGND 
+ VPWR
+ VPWR _0886_ sky130_fd_sc_hd__a22o_1
X_5085_ \gpio_configure[2][10]\ _1486_ net363 _1487_ VGND VGND 
+ VPWR
+ VPWR _0885_ sky130_fd_sc_hd__a22o_1
X_5086_ \gpio_configure[2][9]\ _1486_ net366 _1487_ VGND VGND 
+ VPWR
+ VPWR _0884_ sky130_fd_sc_hd__a22o_1
X_5087_ \gpio_configure[2][8]\ _1486_ net367 _1487_ VGND VGND 
+ VPWR
+ VPWR _0883_ sky130_fd_sc_hd__a22o_1
X_5088_ _1021_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__buf_12
X_5089_ _1488_ _1249_ VGND VGND VPWR VPWR 
+ _1489_
+ sky130_fd_sc_hd__or2_1
X_5090_ _1489_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__buf_2
X_5091_ _1490_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__clkinv_2
X_5092_ \gpio_configure[1][7]\ _1490_ \cdata[7]\ _1491_ VGND VGND 
+ VPWR
+ VPWR _0882_ sky130_fd_sc_hd__a22o_1
X_5093_ \gpio_configure[1][6]\ _1490_ \cdata[6]\ _1491_ VGND VGND 
+ VPWR
+ VPWR _0881_ sky130_fd_sc_hd__a22o_1
X_5094_ \gpio_configure[1][5]\ _1490_ \cdata[5]\ _1491_ VGND VGND 
+ VPWR
+ VPWR _0880_ sky130_fd_sc_hd__a22o_1
X_5095_ \gpio_configure[1][4]\ _1490_ net360 _1491_ VGND VGND 
+ VPWR
+ VPWR _0879_ sky130_fd_sc_hd__a22o_1
X_5096_ \gpio_configure[1][3]\ _1490_ net362 _1491_ VGND VGND 
+ VPWR
+ VPWR _0878_ sky130_fd_sc_hd__a22o_1
X_5097_ \gpio_configure[1][2]\ _1490_ net364 _1491_ VGND VGND 
+ VPWR
+ VPWR _0877_ sky130_fd_sc_hd__a22o_1
X_5098_ \gpio_configure[1][1]\ _1490_ net366 _1491_ VGND VGND 
+ VPWR
+ VPWR _0876_ sky130_fd_sc_hd__a22o_1
X_5099_ \gpio_configure[1][0]\ _1490_ net368 _1491_ VGND VGND 
+ VPWR
+ VPWR _0875_ sky130_fd_sc_hd__a22o_1
X_5100_ _1043_ _1302_ VGND VGND VPWR VPWR 
+ _1492_
+ sky130_fd_sc_hd__or2_1
X_5101_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__clkbuf_2
X_5102_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__inv_2
X_5103_ \gpio_configure[1][12]\ _1493_ net359 _1494_ VGND VGND 
+ VPWR
+ VPWR _0874_ sky130_fd_sc_hd__a22o_1
X_5104_ \gpio_configure[1][11]\ _1493_ net361 _1494_ VGND VGND 
+ VPWR
+ VPWR _0873_ sky130_fd_sc_hd__a22o_1
X_5105_ \gpio_configure[1][10]\ _1493_ net363 _1494_ VGND VGND 
+ VPWR
+ VPWR _0872_ sky130_fd_sc_hd__a22o_1
X_5106_ \gpio_configure[1][9]\ _1493_ net365 _1494_ VGND VGND 
+ VPWR
+ VPWR _0871_ sky130_fd_sc_hd__a22o_1
X_5107_ \gpio_configure[1][8]\ _1493_ net367 _1494_ VGND VGND 
+ VPWR
+ VPWR _0870_ sky130_fd_sc_hd__a22o_1
X_5108_ \wbbd_state[2]\ \wbbd_state[3]\ \wbbd_state[4]\ \wbbd_state[1]\ VGND VGND 
+ VPWR
+ VPWR _1495_ sky130_fd_sc_hd__or4_2
X_5109_ wbbd_sck _1495_ _1080_ _1087_ VGND VGND 
+ VPWR
+ VPWR _0869_ sky130_fd_sc_hd__o211a_2
X_5110_ _1488_ _1353_ VGND VGND VPWR VPWR 
+ _1496_
+ sky130_fd_sc_hd__or2_1
X_5111_ _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__clkbuf_4
X_5112_ _1497_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__inv_2
X_5113_ \gpio_configure[0][7]\ _1497_ \cdata[7]\ _1498_ VGND VGND 
+ VPWR
+ VPWR _0868_ sky130_fd_sc_hd__a22o_1
X_5114_ \gpio_configure[0][6]\ _1497_ \cdata[6]\ _1498_ VGND VGND 
+ VPWR
+ VPWR _0867_ sky130_fd_sc_hd__a22o_1
X_5115_ \gpio_configure[0][5]\ _1497_ \cdata[5]\ _1498_ VGND VGND 
+ VPWR
+ VPWR _0866_ sky130_fd_sc_hd__a22o_1
X_5116_ \gpio_configure[0][4]\ _1497_ net359 _1498_ VGND VGND 
+ VPWR
+ VPWR _0865_ sky130_fd_sc_hd__a22o_1
X_5117_ \gpio_configure[0][3]\ _1497_ net361 _1498_ VGND VGND 
+ VPWR
+ VPWR _0864_ sky130_fd_sc_hd__a22o_1
X_5118_ \gpio_configure[0][2]\ _1497_ net363 _1498_ VGND VGND 
+ VPWR
+ VPWR _0863_ sky130_fd_sc_hd__a22o_1
X_5119_ \gpio_configure[0][1]\ _1497_ net365 _1498_ VGND VGND 
+ VPWR
+ VPWR _0862_ sky130_fd_sc_hd__a22o_1
X_5120_ \gpio_configure[0][0]\ _1497_ net367 _1498_ VGND VGND 
+ VPWR
+ VPWR _0861_ sky130_fd_sc_hd__a22o_1
X_5121_ _1043_ _1275_ VGND VGND VPWR VPWR 
+ _1499_
+ sky130_fd_sc_hd__or2_1
X_5122_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__clkbuf_2
X_5123_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__inv_2
X_5124_ \gpio_configure[0][12]\ _1500_ net359 _1501_ VGND VGND 
+ VPWR
+ VPWR _0860_ sky130_fd_sc_hd__a22o_1
X_5125_ \gpio_configure[0][11]\ _1500_ net361 _1501_ VGND VGND 
+ VPWR
+ VPWR _0859_ sky130_fd_sc_hd__a22o_1
X_5126_ \gpio_configure[0][10]\ _1500_ net363 _1501_ VGND VGND 
+ VPWR
+ VPWR _0858_ sky130_fd_sc_hd__a22o_1
X_5127_ \gpio_configure[0][9]\ _1500_ net365 _1501_ VGND VGND 
+ VPWR
+ VPWR _0857_ sky130_fd_sc_hd__a22o_1
X_5128_ \gpio_configure[0][8]\ _1500_ net367 _1501_ VGND VGND 
+ VPWR
+ VPWR _0856_ sky130_fd_sc_hd__a22o_1
X_5129_ _1449_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__clkbuf_1
X_5130_ _1502_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_5131_ \hkspi.state[0]\ _1423_ \hkspi.pre_pass_thru_mgmt\ \hkspi.pass_thru_mgmt_delay\ _1424_ VGND 
+ VGND
+ VPWR VPWR _0855_ sky130_fd_sc_hd__a32o_1
X_5132_ _1125_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__inv_8
X_5133_ _1021_ _0079_ VGND VGND VPWR VPWR 
+ _1503_
+ sky130_fd_sc_hd__or2_4
X_5134_ _1177_ _1503_ VGND VGND VPWR VPWR 
+ _1504_
+ sky130_fd_sc_hd__or2_1
X_5135_ _1504_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__clkbuf_4
X_5136_ _1505_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__inv_2
X_5137_ \mgmt_gpio_data_buf[7]\ _1505_ \cdata[7]\ _1506_ VGND VGND 
+ VPWR
+ VPWR _0854_ sky130_fd_sc_hd__a22o_1
X_5138_ \mgmt_gpio_data_buf[6]\ _1505_ \cdata[6]\ _1506_ VGND VGND 
+ VPWR
+ VPWR _0853_ sky130_fd_sc_hd__a22o_1
X_5139_ \mgmt_gpio_data_buf[5]\ _1505_ \cdata[5]\ _1506_ VGND VGND 
+ VPWR
+ VPWR _0852_ sky130_fd_sc_hd__a22o_1
X_5140_ \mgmt_gpio_data_buf[4]\ _1505_ net360 _1506_ VGND VGND 
+ VPWR
+ VPWR _0851_ sky130_fd_sc_hd__a22o_1
X_5141_ \mgmt_gpio_data_buf[3]\ _1505_ net362 _1506_ VGND VGND 
+ VPWR
+ VPWR _0850_ sky130_fd_sc_hd__a22o_1
X_5142_ \mgmt_gpio_data_buf[2]\ _1505_ net364 _1506_ VGND VGND 
+ VPWR
+ VPWR _0849_ sky130_fd_sc_hd__a22o_1
X_5143_ \mgmt_gpio_data_buf[1]\ _1505_ net366 _1506_ VGND VGND 
+ VPWR
+ VPWR _0848_ sky130_fd_sc_hd__a22o_1
X_5144_ \mgmt_gpio_data_buf[0]\ _1505_ net368 _1506_ VGND VGND 
+ VPWR
+ VPWR _0847_ sky130_fd_sc_hd__a22o_1
X_5145_ _1218_ _1503_ VGND VGND VPWR VPWR 
+ _1507_
+ sky130_fd_sc_hd__or2_1
X_5146_ _1507_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__clkbuf_4
X_5147_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__inv_2
X_5148_ \mgmt_gpio_data_buf[15]\ _1508_ \cdata[7]\ _1509_ VGND VGND 
+ VPWR
+ VPWR _0846_ sky130_fd_sc_hd__a22o_1
X_5149_ \mgmt_gpio_data_buf[14]\ _1508_ \cdata[6]\ _1509_ VGND VGND 
+ VPWR
+ VPWR _0845_ sky130_fd_sc_hd__a22o_1
X_5150_ \mgmt_gpio_data_buf[13]\ _1508_ \cdata[5]\ _1509_ VGND VGND 
+ VPWR
+ VPWR _0844_ sky130_fd_sc_hd__a22o_1
X_5151_ \mgmt_gpio_data_buf[12]\ _1508_ net360 _1509_ VGND VGND 
+ VPWR
+ VPWR _0843_ sky130_fd_sc_hd__a22o_1
X_5152_ \mgmt_gpio_data_buf[11]\ _1508_ net362 _1509_ VGND VGND 
+ VPWR
+ VPWR _0842_ sky130_fd_sc_hd__a22o_1
X_5153_ \mgmt_gpio_data_buf[10]\ _1508_ net364 _1509_ VGND VGND 
+ VPWR
+ VPWR _0841_ sky130_fd_sc_hd__a22o_1
X_5154_ \mgmt_gpio_data_buf[9]\ _1508_ net366 _1509_ VGND VGND 
+ VPWR
+ VPWR _0840_ sky130_fd_sc_hd__a22o_1
X_5155_ \mgmt_gpio_data_buf[8]\ _1508_ net368 _1509_ VGND VGND 
+ VPWR
+ VPWR _0839_ sky130_fd_sc_hd__a22o_1
X_5156_ _1235_ _1503_ VGND VGND VPWR VPWR 
+ _1510_
+ sky130_fd_sc_hd__or2_1
X_5157_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__clkbuf_4
X_5158_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__inv_2
X_5159_ \mgmt_gpio_data_buf[23]\ _1511_ \cdata[7]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0838_ sky130_fd_sc_hd__a22o_1
X_5160_ \mgmt_gpio_data_buf[22]\ _1511_ \cdata[6]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0837_ sky130_fd_sc_hd__a22o_1
X_5161_ \mgmt_gpio_data_buf[21]\ _1511_ \cdata[5]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0836_ sky130_fd_sc_hd__a22o_1
X_5162_ \mgmt_gpio_data_buf[20]\ _1511_ net360 _1512_ VGND VGND 
+ VPWR
+ VPWR _0835_ sky130_fd_sc_hd__a22o_1
X_5163_ \mgmt_gpio_data_buf[19]\ _1511_ \cdata[3]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0834_ sky130_fd_sc_hd__a22o_1
X_5164_ \mgmt_gpio_data_buf[18]\ _1511_ \cdata[2]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0833_ sky130_fd_sc_hd__a22o_1
X_5165_ \mgmt_gpio_data_buf[17]\ _1511_ \cdata[1]\ _1512_ VGND VGND 
+ VPWR
+ VPWR _0832_ sky130_fd_sc_hd__a22o_1
X_5166_ \mgmt_gpio_data_buf[16]\ _1511_ net368 _1512_ VGND VGND 
+ VPWR
+ VPWR _0831_ sky130_fd_sc_hd__a22o_1
X_5167_ _1488_ _1262_ VGND VGND VPWR VPWR 
+ _1513_
+ sky130_fd_sc_hd__or2_1
X_5168_ _1513_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__clkbuf_4
X_5169_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__inv_2
X_5170_ \mgmt_gpio_data[31]\ _1514_ \cdata[7]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0830_ sky130_fd_sc_hd__a22o_1
X_5171_ \mgmt_gpio_data[30]\ _1514_ \cdata[6]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0829_ sky130_fd_sc_hd__a22o_1
X_5172_ \mgmt_gpio_data[29]\ _1514_ \cdata[5]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0828_ sky130_fd_sc_hd__a22o_1
X_5173_ \mgmt_gpio_data[28]\ _1514_ net360 _1515_ VGND VGND 
+ VPWR
+ VPWR _0827_ sky130_fd_sc_hd__a22o_1
X_5174_ \mgmt_gpio_data[27]\ _1514_ \cdata[3]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0826_ sky130_fd_sc_hd__a22o_1
X_5175_ \mgmt_gpio_data[26]\ _1514_ \cdata[2]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0825_ sky130_fd_sc_hd__a22o_1
X_5176_ \mgmt_gpio_data[25]\ _1514_ \cdata[1]\ _1515_ VGND VGND 
+ VPWR
+ VPWR _0824_ sky130_fd_sc_hd__a22o_1
X_5177_ \mgmt_gpio_data[24]\ _1514_ net368 _1515_ VGND VGND 
+ VPWR
+ VPWR _0823_ sky130_fd_sc_hd__a22o_1
X_5178_ _1023_ _1158_ VGND VGND VPWR VPWR 
+ _1516_
+ sky130_fd_sc_hd__or2_2
X_5179_ _1516_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__buf_2
X_5180_ _1517_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__clkinv_2
X_5181_ \mgmt_gpio_data[37]\ _1517_ \cdata[5]\ _1518_ VGND VGND 
+ VPWR
+ VPWR _0822_ sky130_fd_sc_hd__a22o_1
X_5182_ \mgmt_gpio_data[36]\ _1517_ net360 _1518_ VGND VGND 
+ VPWR
+ VPWR _0821_ sky130_fd_sc_hd__a22o_1
X_5183_ \mgmt_gpio_data[35]\ _1517_ \cdata[3]\ _1518_ VGND VGND 
+ VPWR
+ VPWR _0820_ sky130_fd_sc_hd__a22o_1
X_5184_ \mgmt_gpio_data[34]\ _1517_ \cdata[2]\ _1518_ VGND VGND 
+ VPWR
+ VPWR _0819_ sky130_fd_sc_hd__a22o_1
X_5185_ \mgmt_gpio_data[33]\ _1517_ \cdata[1]\ _1518_ VGND VGND 
+ VPWR
+ VPWR _0818_ sky130_fd_sc_hd__a22o_1
X_5186_ \mgmt_gpio_data[32]\ _1517_ net368 _1518_ VGND VGND 
+ VPWR
+ VPWR _0817_ sky130_fd_sc_hd__a22o_1
X_5187_ \wbbd_state[0]\ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__inv_2
X_5188_ wbbd_busy _1519_ _1495_ _1088_ VGND VGND 
+ VPWR
+ VPWR _0816_ sky130_fd_sc_hd__a211o_1
X_5189_ _1449_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__clkbuf_1
X_5190_ _1520_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
X_5191_ \hkspi.state[4]\ _1466_ \hkspi.pass_thru_mgmt\ VGND VGND VPWR 
+ VPWR
+ _0815_ sky130_fd_sc_hd__a21o_1
X_5192_ _1262_ _1177_ _1043_ _0086_ VGND VGND 
+ VPWR
+ VPWR _1521_ sky130_fd_sc_hd__a211o_4
X_5193_ _1521_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__inv_2
X_5194_ \mgmt_gpio_data[7]\ _1522_ _0199_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0814_ sky130_fd_sc_hd__o22a_1
X_5195_ \mgmt_gpio_data[6]\ _1522_ _0198_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0813_ sky130_fd_sc_hd__o22a_1
X_5196_ \mgmt_gpio_data[5]\ _1522_ _0197_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0812_ sky130_fd_sc_hd__o22a_1
X_5197_ \mgmt_gpio_data[4]\ _1522_ _0196_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0811_ sky130_fd_sc_hd__o22a_1
X_5198_ \mgmt_gpio_data[3]\ _1522_ _0195_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0810_ sky130_fd_sc_hd__o22a_1
X_5199_ \mgmt_gpio_data[2]\ _1522_ _0194_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0809_ sky130_fd_sc_hd__o22a_1
X_5200_ \mgmt_gpio_data[1]\ _1522_ _0193_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0808_ sky130_fd_sc_hd__o22a_1
X_5201_ \mgmt_gpio_data[0]\ _1522_ _0192_ _1521_ VGND VGND 
+ VPWR
+ VPWR _0807_ sky130_fd_sc_hd__o22a_1
X_5202_ _1218_ _1262_ _1043_ _0084_ VGND VGND 
+ VPWR
+ VPWR _1523_ sky130_fd_sc_hd__a211o_4
X_5203_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__inv_2
X_5204_ \mgmt_gpio_data[15]\ _1524_ _0207_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0806_ sky130_fd_sc_hd__o22a_1
X_5205_ \mgmt_gpio_data[14]\ _1524_ _0206_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0805_ sky130_fd_sc_hd__o22a_1
X_5206_ \mgmt_gpio_data[13]\ _1524_ _0205_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0804_ sky130_fd_sc_hd__o22a_1
X_5207_ \mgmt_gpio_data[12]\ _1524_ _0204_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0803_ sky130_fd_sc_hd__o22a_1
X_5208_ \mgmt_gpio_data[11]\ _1524_ _0203_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0802_ sky130_fd_sc_hd__o22a_1
X_5209_ \mgmt_gpio_data[10]\ _1524_ _0202_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0801_ sky130_fd_sc_hd__o22a_1
X_5210_ \mgmt_gpio_data[9]\ _1524_ _0201_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0800_ sky130_fd_sc_hd__o22a_1
X_5211_ \mgmt_gpio_data[8]\ _1524_ _0200_ _1523_ VGND VGND 
+ VPWR
+ VPWR _0799_ sky130_fd_sc_hd__o22a_1
X_5212_ _1449_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__clkbuf_1
X_5213_ _1525_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
X_5214_ _0154_ _1466_ VGND VGND VPWR VPWR 
+ _1526_
+ sky130_fd_sc_hd__nor2_1
X_5215_ \hkspi.state[0]\ _1419_ VGND VGND VPWR VPWR 
+ _1527_
+ sky130_fd_sc_hd__nor2_1
X_5216_ \hkspi.rdstb\ _1526_ _1466_ _1527_ VGND VGND 
+ VPWR
+ VPWR _0798_ sky130_fd_sc_hd__o22a_1
X_5217_ _1235_ _1262_ _1043_ _0082_ VGND VGND 
+ VPWR
+ VPWR _1528_ sky130_fd_sc_hd__a211o_4
X_5218_ _1528_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__inv_2
X_5219_ \mgmt_gpio_data[23]\ _1529_ _0215_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0797_ sky130_fd_sc_hd__o22a_1
X_5220_ \mgmt_gpio_data[22]\ _1529_ _0214_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0796_ sky130_fd_sc_hd__o22a_1
X_5221_ \mgmt_gpio_data[21]\ _1529_ _0213_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0795_ sky130_fd_sc_hd__o22a_1
X_5222_ \mgmt_gpio_data[20]\ _1529_ _0212_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0794_ sky130_fd_sc_hd__o22a_1
X_5223_ \mgmt_gpio_data[19]\ _1529_ _0211_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0793_ sky130_fd_sc_hd__o22a_1
X_5224_ \mgmt_gpio_data[18]\ _1529_ _0210_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0792_ sky130_fd_sc_hd__o22a_1
X_5225_ \mgmt_gpio_data[17]\ _1529_ _0209_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0791_ sky130_fd_sc_hd__o22a_1
X_5226_ \mgmt_gpio_data[16]\ _1529_ _0208_ _1528_ VGND VGND 
+ VPWR
+ VPWR _0790_ sky130_fd_sc_hd__o22a_1
X_5227_ _1043_ _1304_ VGND VGND VPWR VPWR 
+ _1530_
+ sky130_fd_sc_hd__or2_1
X_5228_ net365 irq_2_inputsrc _1530_ VGND VGND VPWR 
+ VPWR
+ _1531_ sky130_fd_sc_hd__mux2_1
X_5229_ _1531_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__clkbuf_1
X_5230_ net367 irq_1_inputsrc _1530_ VGND VGND VPWR 
+ VPWR
+ _1532_ sky130_fd_sc_hd__mux2_1
X_5231_ _1532_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__clkbuf_1
X_5232_ _1043_ _1315_ VGND VGND VPWR VPWR 
+ _1533_
+ sky130_fd_sc_hd__or2_1
X_5233_ _1533_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__clkbuf_2
X_5234_ _1534_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__inv_2
X_5235_ \gpio_configure[27][12]\ _1534_ net359 _1535_ VGND VGND 
+ VPWR
+ VPWR _0787_ sky130_fd_sc_hd__a22o_1
X_5236_ \gpio_configure[27][11]\ _1534_ net361 _1535_ VGND VGND 
+ VPWR
+ VPWR _0786_ sky130_fd_sc_hd__a22o_1
X_5237_ \gpio_configure[27][10]\ _1534_ net363 _1535_ VGND VGND 
+ VPWR
+ VPWR _0785_ sky130_fd_sc_hd__a22o_1
X_5238_ \gpio_configure[27][9]\ _1534_ net365 _1535_ VGND VGND 
+ VPWR
+ VPWR _0784_ sky130_fd_sc_hd__a22o_1
X_5239_ \gpio_configure[27][8]\ _1534_ net367 _1535_ VGND VGND 
+ VPWR
+ VPWR _0783_ sky130_fd_sc_hd__a22o_1
X_5240_ _1488_ _1273_ VGND VGND VPWR VPWR 
+ _1536_
+ sky130_fd_sc_hd__or2_1
X_5241_ _1536_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__clkbuf_4
X_5242_ _1537_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__inv_2
X_5243_ \gpio_configure[27][7]\ _1537_ \cdata[7]\ _1538_ VGND VGND 
+ VPWR
+ VPWR _0782_ sky130_fd_sc_hd__a22o_1
X_5244_ \gpio_configure[27][6]\ _1537_ \cdata[6]\ _1538_ VGND VGND 
+ VPWR
+ VPWR _0781_ sky130_fd_sc_hd__a22o_1
X_5245_ \gpio_configure[27][5]\ _1537_ \cdata[5]\ _1538_ VGND VGND 
+ VPWR
+ VPWR _0780_ sky130_fd_sc_hd__a22o_1
X_5246_ \gpio_configure[27][4]\ _1537_ net359 _1538_ VGND VGND 
+ VPWR
+ VPWR _0779_ sky130_fd_sc_hd__a22o_1
X_5247_ \gpio_configure[27][3]\ _1537_ net361 _1538_ VGND VGND 
+ VPWR
+ VPWR _0778_ sky130_fd_sc_hd__a22o_1
X_5248_ \gpio_configure[27][2]\ _1537_ net363 _1538_ VGND VGND 
+ VPWR
+ VPWR _0777_ sky130_fd_sc_hd__a22o_1
X_5249_ \gpio_configure[27][1]\ _1537_ net365 _1538_ VGND VGND 
+ VPWR
+ VPWR _0776_ sky130_fd_sc_hd__a22o_1
X_5250_ \gpio_configure[27][0]\ _1537_ net367 _1538_ VGND VGND 
+ VPWR
+ VPWR _0775_ sky130_fd_sc_hd__a22o_1
X_5251_ _1043_ _1288_ VGND VGND VPWR VPWR 
+ _1539_
+ sky130_fd_sc_hd__or2_1
X_5252_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__clkbuf_2
X_5253_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__inv_2
X_5254_ \gpio_configure[25][12]\ _1540_ net359 _1541_ VGND VGND 
+ VPWR
+ VPWR _0774_ sky130_fd_sc_hd__a22o_1
X_5255_ \gpio_configure[25][11]\ _1540_ net361 _1541_ VGND VGND 
+ VPWR
+ VPWR _0773_ sky130_fd_sc_hd__a22o_1
X_5256_ \gpio_configure[25][10]\ _1540_ net363 _1541_ VGND VGND 
+ VPWR
+ VPWR _0772_ sky130_fd_sc_hd__a22o_1
X_5257_ \gpio_configure[25][9]\ _1540_ net365 _1541_ VGND VGND 
+ VPWR
+ VPWR _0771_ sky130_fd_sc_hd__a22o_1
X_5258_ \gpio_configure[25][8]\ _1540_ net367 _1541_ VGND VGND 
+ VPWR
+ VPWR _0770_ sky130_fd_sc_hd__a22o_1
X_5259_ _1043_ _1361_ VGND VGND VPWR VPWR 
+ _1542_
+ sky130_fd_sc_hd__or2_1
X_5260_ _1542_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__clkbuf_2
X_5261_ _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__inv_2
X_5262_ \gpio_configure[28][12]\ _1543_ net359 _1544_ VGND VGND 
+ VPWR
+ VPWR _0769_ sky130_fd_sc_hd__a22o_1
X_5263_ \gpio_configure[28][11]\ _1543_ net361 _1544_ VGND VGND 
+ VPWR
+ VPWR _0768_ sky130_fd_sc_hd__a22o_1
X_5264_ \gpio_configure[28][10]\ _1543_ net363 _1544_ VGND VGND 
+ VPWR
+ VPWR _0767_ sky130_fd_sc_hd__a22o_1
X_5265_ \gpio_configure[28][9]\ _1543_ net365 _1544_ VGND VGND 
+ VPWR
+ VPWR _0766_ sky130_fd_sc_hd__a22o_1
X_5266_ \gpio_configure[28][8]\ _1543_ net367 _1544_ VGND VGND 
+ VPWR
+ VPWR _0765_ sky130_fd_sc_hd__a22o_1
X_5267_ _1488_ _1325_ VGND VGND VPWR VPWR 
+ _1545_
+ sky130_fd_sc_hd__or2_1
X_5268_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__buf_2
X_5269_ _1546_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__clkinv_2
X_5270_ \gpio_configure[24][7]\ _1546_ \cdata[7]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0764_ sky130_fd_sc_hd__a22o_1
X_5271_ \gpio_configure[24][6]\ _1546_ \cdata[6]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0763_ sky130_fd_sc_hd__a22o_1
X_5272_ \gpio_configure[24][5]\ _1546_ \cdata[5]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0762_ sky130_fd_sc_hd__a22o_1
X_5273_ \gpio_configure[24][4]\ _1546_ \cdata[4]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0761_ sky130_fd_sc_hd__a22o_1
X_5274_ \gpio_configure[24][3]\ _1546_ net362 _1547_ VGND VGND 
+ VPWR
+ VPWR _0760_ sky130_fd_sc_hd__a22o_1
X_5275_ \gpio_configure[24][2]\ _1546_ \cdata[2]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0759_ sky130_fd_sc_hd__a22o_1
X_5276_ \gpio_configure[24][1]\ _1546_ net366 _1547_ VGND VGND 
+ VPWR
+ VPWR _0758_ sky130_fd_sc_hd__a22o_1
X_5277_ \gpio_configure[24][0]\ _1546_ \cdata[0]\ _1547_ VGND VGND 
+ VPWR
+ VPWR _0757_ sky130_fd_sc_hd__a22o_1
X_5278_ _1488_ _1388_ VGND VGND VPWR VPWR 
+ _1548_
+ sky130_fd_sc_hd__or2_1
X_5279_ _1548_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__clkbuf_4
X_5280_ _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__inv_2
X_5281_ \gpio_configure[28][7]\ _1549_ \cdata[7]\ _1550_ VGND VGND 
+ VPWR
+ VPWR _0756_ sky130_fd_sc_hd__a22o_1
X_5282_ \gpio_configure[28][6]\ _1549_ \cdata[6]\ _1550_ VGND VGND 
+ VPWR
+ VPWR _0755_ sky130_fd_sc_hd__a22o_1
X_5283_ \gpio_configure[28][5]\ _1549_ \cdata[5]\ _1550_ VGND VGND 
+ VPWR
+ VPWR _0754_ sky130_fd_sc_hd__a22o_1
X_5284_ \gpio_configure[28][4]\ _1549_ net360 _1550_ VGND VGND 
+ VPWR
+ VPWR _0753_ sky130_fd_sc_hd__a22o_1
X_5285_ \gpio_configure[28][3]\ _1549_ \cdata[3]\ _1550_ VGND VGND 
+ VPWR
+ VPWR _0752_ sky130_fd_sc_hd__a22o_1
X_5286_ \gpio_configure[28][2]\ _1549_ net364 _1550_ VGND VGND 
+ VPWR
+ VPWR _0751_ sky130_fd_sc_hd__a22o_1
X_5287_ \gpio_configure[28][1]\ _1549_ \cdata[1]\ _1550_ VGND VGND 
+ VPWR
+ VPWR _0750_ sky130_fd_sc_hd__a22o_1
X_5288_ \gpio_configure[28][0]\ _1549_ net368 _1550_ VGND VGND 
+ VPWR
+ VPWR _0749_ sky130_fd_sc_hd__a22o_1
X_5289_ _1022_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__clkbuf_16
X_5290_ _1551_ _1282_ VGND VGND VPWR VPWR 
+ _1552_
+ sky130_fd_sc_hd__or2_1
X_5291_ _1552_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__clkbuf_2
X_5292_ _1553_ VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__inv_2
X_5293_ \gpio_configure[24][12]\ _1553_ net359 _1554_ VGND VGND 
+ VPWR
+ VPWR _0748_ sky130_fd_sc_hd__a22o_1
X_5294_ \gpio_configure[24][11]\ _1553_ net361 _1554_ VGND VGND 
+ VPWR
+ VPWR _0747_ sky130_fd_sc_hd__a22o_1
X_5295_ \gpio_configure[24][10]\ _1553_ net363 _1554_ VGND VGND 
+ VPWR
+ VPWR _0746_ sky130_fd_sc_hd__a22o_1
X_5296_ \gpio_configure[24][9]\ _1553_ net365 _1554_ VGND VGND 
+ VPWR
+ VPWR _0745_ sky130_fd_sc_hd__a22o_1
X_5297_ \gpio_configure[24][8]\ _1553_ net367 _1554_ VGND VGND 
+ VPWR
+ VPWR _0744_ sky130_fd_sc_hd__a22o_1
X_5298_ _1551_ _1366_ VGND VGND VPWR VPWR 
+ _1555_
+ sky130_fd_sc_hd__or2_1
X_5299_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__clkbuf_2
X_5300_ _1556_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__inv_2
X_5301_ \gpio_configure[29][12]\ _1556_ net359 _1557_ VGND VGND 
+ VPWR
+ VPWR _0743_ sky130_fd_sc_hd__a22o_1
X_5302_ \gpio_configure[29][11]\ _1556_ net361 _1557_ VGND VGND 
+ VPWR
+ VPWR _0742_ sky130_fd_sc_hd__a22o_1
X_5303_ \gpio_configure[29][10]\ _1556_ net363 _1557_ VGND VGND 
+ VPWR
+ VPWR _0741_ sky130_fd_sc_hd__a22o_1
X_5304_ \gpio_configure[29][9]\ _1556_ net365 _1557_ VGND VGND 
+ VPWR
+ VPWR _0740_ sky130_fd_sc_hd__a22o_1
X_5305_ \gpio_configure[29][8]\ _1556_ net367 _1557_ VGND VGND 
+ VPWR
+ VPWR _0739_ sky130_fd_sc_hd__a22o_1
X_5306_ _1488_ _1404_ VGND VGND VPWR VPWR 
+ _1558_
+ sky130_fd_sc_hd__or2_1
X_5307_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__clkbuf_4
X_5308_ _1559_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__inv_2
X_5309_ \gpio_configure[23][7]\ _1559_ \cdata[7]\ _1560_ VGND VGND 
+ VPWR
+ VPWR _0738_ sky130_fd_sc_hd__a22o_1
X_5310_ \gpio_configure[23][6]\ _1559_ \cdata[6]\ _1560_ VGND VGND 
+ VPWR
+ VPWR _0737_ sky130_fd_sc_hd__a22o_1
X_5311_ \gpio_configure[23][5]\ _1559_ \cdata[5]\ _1560_ VGND VGND 
+ VPWR
+ VPWR _0736_ sky130_fd_sc_hd__a22o_1
X_5312_ \gpio_configure[23][4]\ _1559_ net360 _1560_ VGND VGND 
+ VPWR
+ VPWR _0735_ sky130_fd_sc_hd__a22o_1
X_5313_ \gpio_configure[23][3]\ _1559_ \cdata[3]\ _1560_ VGND VGND 
+ VPWR
+ VPWR _0734_ sky130_fd_sc_hd__a22o_1
X_5314_ \gpio_configure[23][2]\ _1559_ net364 _1560_ VGND VGND 
+ VPWR
+ VPWR _0733_ sky130_fd_sc_hd__a22o_1
X_5315_ \gpio_configure[23][1]\ _1559_ \cdata[1]\ _1560_ VGND VGND 
+ VPWR
+ VPWR _0732_ sky130_fd_sc_hd__a22o_1
X_5316_ \gpio_configure[23][0]\ _1559_ net368 _1560_ VGND VGND 
+ VPWR
+ VPWR _0731_ sky130_fd_sc_hd__a22o_1
X_5317_ _1488_ _1334_ VGND VGND VPWR VPWR 
+ _1561_
+ sky130_fd_sc_hd__or2_1
X_5318_ _1561_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__clkbuf_4
X_5319_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__inv_2
X_5320_ \gpio_configure[29][7]\ _1562_ \cdata[7]\ _1563_ VGND VGND 
+ VPWR
+ VPWR _0730_ sky130_fd_sc_hd__a22o_1
X_5321_ \gpio_configure[29][6]\ _1562_ \cdata[6]\ _1563_ VGND VGND 
+ VPWR
+ VPWR _0729_ sky130_fd_sc_hd__a22o_1
X_5322_ \gpio_configure[29][5]\ _1562_ \cdata[5]\ _1563_ VGND VGND 
+ VPWR
+ VPWR _0728_ sky130_fd_sc_hd__a22o_1
X_5323_ \gpio_configure[29][4]\ _1562_ net360 _1563_ VGND VGND 
+ VPWR
+ VPWR _0727_ sky130_fd_sc_hd__a22o_1
X_5324_ \gpio_configure[29][3]\ _1562_ net362 _1563_ VGND VGND 
+ VPWR
+ VPWR _0726_ sky130_fd_sc_hd__a22o_1
X_5325_ \gpio_configure[29][2]\ _1562_ \cdata[2]\ _1563_ VGND VGND 
+ VPWR
+ VPWR _0725_ sky130_fd_sc_hd__a22o_1
X_5326_ \gpio_configure[29][1]\ _1562_ net366 _1563_ VGND VGND 
+ VPWR
+ VPWR _0724_ sky130_fd_sc_hd__a22o_1
X_5327_ \gpio_configure[29][0]\ _1562_ \cdata[0]\ _1563_ VGND VGND 
+ VPWR
+ VPWR _0723_ sky130_fd_sc_hd__a22o_1
X_5328_ _1551_ _1408_ VGND VGND VPWR VPWR 
+ _1564_
+ sky130_fd_sc_hd__or2_1
X_5329_ _1564_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__clkbuf_2
X_5330_ _1565_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__inv_2
X_5331_ \gpio_configure[23][12]\ _1565_ net359 _1566_ VGND VGND 
+ VPWR
+ VPWR _0722_ sky130_fd_sc_hd__a22o_1
X_5332_ \gpio_configure[23][11]\ _1565_ net361 _1566_ VGND VGND 
+ VPWR
+ VPWR _0721_ sky130_fd_sc_hd__a22o_1
X_5333_ \gpio_configure[23][10]\ _1565_ net363 _1566_ VGND VGND 
+ VPWR
+ VPWR _0720_ sky130_fd_sc_hd__a22o_1
X_5334_ \gpio_configure[23][9]\ _1565_ net365 _1566_ VGND VGND 
+ VPWR
+ VPWR _0719_ sky130_fd_sc_hd__a22o_1
X_5335_ \gpio_configure[23][8]\ _1565_ net367 _1566_ VGND VGND 
+ VPWR
+ VPWR _0718_ sky130_fd_sc_hd__a22o_1
X_5336_ _1551_ _1344_ VGND VGND VPWR VPWR 
+ _1567_
+ sky130_fd_sc_hd__or2_1
X_5337_ _1567_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__clkbuf_2
X_5338_ _1568_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__inv_2
X_5339_ \gpio_configure[30][12]\ _1568_ net359 _1569_ VGND VGND 
+ VPWR
+ VPWR _0717_ sky130_fd_sc_hd__a22o_1
X_5340_ \gpio_configure[30][11]\ _1568_ net361 _1569_ VGND VGND 
+ VPWR
+ VPWR _0716_ sky130_fd_sc_hd__a22o_1
X_5341_ \gpio_configure[30][10]\ _1568_ net363 _1569_ VGND VGND 
+ VPWR
+ VPWR _0715_ sky130_fd_sc_hd__a22o_1
X_5342_ \gpio_configure[30][9]\ _1568_ net365 _1569_ VGND VGND 
+ VPWR
+ VPWR _0714_ sky130_fd_sc_hd__a22o_1
X_5343_ \gpio_configure[30][8]\ _1568_ net367 _1569_ VGND VGND 
+ VPWR
+ VPWR _0713_ sky130_fd_sc_hd__a22o_1
X_5344_ _1488_ _1375_ VGND VGND VPWR VPWR 
+ _1570_
+ sky130_fd_sc_hd__or2_1
X_5345_ _1570_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__clkbuf_4
X_5346_ _1571_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__inv_2
X_5347_ \gpio_configure[22][7]\ _1571_ \cdata[7]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0712_ sky130_fd_sc_hd__a22o_1
X_5348_ \gpio_configure[22][6]\ _1571_ \cdata[6]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0711_ sky130_fd_sc_hd__a22o_1
X_5349_ \gpio_configure[22][5]\ _1571_ \cdata[5]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0710_ sky130_fd_sc_hd__a22o_1
X_5350_ \gpio_configure[22][4]\ _1571_ net360 _1572_ VGND VGND 
+ VPWR
+ VPWR _0709_ sky130_fd_sc_hd__a22o_1
X_5351_ \gpio_configure[22][3]\ _1571_ \cdata[3]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0708_ sky130_fd_sc_hd__a22o_1
X_5352_ \gpio_configure[22][2]\ _1571_ \cdata[2]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0707_ sky130_fd_sc_hd__a22o_1
X_5353_ \gpio_configure[22][1]\ _1571_ \cdata[1]\ _1572_ VGND VGND 
+ VPWR
+ VPWR _0706_ sky130_fd_sc_hd__a22o_1
X_5354_ \gpio_configure[22][0]\ _1571_ net368 _1572_ VGND VGND 
+ VPWR
+ VPWR _0705_ sky130_fd_sc_hd__a22o_1
X_5355_ _1488_ _1329_ VGND VGND VPWR VPWR 
+ _1573_
+ sky130_fd_sc_hd__or2_1
X_5356_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__clkbuf_4
X_5357_ _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__clkinv_2
X_5358_ \gpio_configure[30][7]\ _1574_ \cdata[7]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0704_ sky130_fd_sc_hd__a22o_1
X_5359_ \gpio_configure[30][6]\ _1574_ \cdata[6]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0703_ sky130_fd_sc_hd__a22o_1
X_5360_ \gpio_configure[30][5]\ _1574_ \cdata[5]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0702_ sky130_fd_sc_hd__a22o_1
X_5361_ \gpio_configure[30][4]\ _1574_ net360 _1575_ VGND VGND 
+ VPWR
+ VPWR _0701_ sky130_fd_sc_hd__a22o_1
X_5362_ \gpio_configure[30][3]\ _1574_ \cdata[3]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0700_ sky130_fd_sc_hd__a22o_1
X_5363_ \gpio_configure[30][2]\ _1574_ \cdata[2]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0699_ sky130_fd_sc_hd__a22o_1
X_5364_ \gpio_configure[30][1]\ _1574_ \cdata[1]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0698_ sky130_fd_sc_hd__a22o_1
X_5365_ \gpio_configure[30][0]\ _1574_ \cdata[0]\ _1575_ VGND VGND 
+ VPWR
+ VPWR _0697_ sky130_fd_sc_hd__a22o_1
X_5366_ _1551_ _1402_ VGND VGND VPWR VPWR 
+ _1576_
+ sky130_fd_sc_hd__or2_1
X_5367_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__clkbuf_2
X_5368_ _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__inv_2
X_5369_ \gpio_configure[22][12]\ _1577_ net359 _1578_ VGND VGND 
+ VPWR
+ VPWR _0696_ sky130_fd_sc_hd__a22o_1
X_5370_ \gpio_configure[22][11]\ _1577_ net361 _1578_ VGND VGND 
+ VPWR
+ VPWR _0695_ sky130_fd_sc_hd__a22o_1
X_5371_ \gpio_configure[22][10]\ _1577_ net363 _1578_ VGND VGND 
+ VPWR
+ VPWR _0694_ sky130_fd_sc_hd__a22o_1
X_5372_ \gpio_configure[22][9]\ _1577_ net365 _1578_ VGND VGND 
+ VPWR
+ VPWR _0693_ sky130_fd_sc_hd__a22o_1
X_5373_ \gpio_configure[22][8]\ _1577_ net367 _1578_ VGND VGND 
+ VPWR
+ VPWR _0692_ sky130_fd_sc_hd__a22o_1
X_5374_ _1551_ _1337_ VGND VGND VPWR VPWR 
+ _1579_
+ sky130_fd_sc_hd__or2_1
X_5375_ _1579_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__clkbuf_2
X_5376_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__inv_2
X_5377_ \gpio_configure[31][12]\ _1580_ \cdata[4]\ _1581_ VGND VGND 
+ VPWR
+ VPWR _0691_ sky130_fd_sc_hd__a22o_1
X_5378_ \gpio_configure[31][11]\ _1580_ \cdata[3]\ _1581_ VGND VGND 
+ VPWR
+ VPWR _0690_ sky130_fd_sc_hd__a22o_1
X_5379_ \gpio_configure[31][10]\ _1580_ \cdata[2]\ _1581_ VGND VGND 
+ VPWR
+ VPWR _0689_ sky130_fd_sc_hd__a22o_1
X_5380_ \gpio_configure[31][9]\ _1580_ net366 _1581_ VGND VGND 
+ VPWR
+ VPWR _0688_ sky130_fd_sc_hd__a22o_1
X_5381_ \gpio_configure[31][8]\ _1580_ \cdata[0]\ _1581_ VGND VGND 
+ VPWR
+ VPWR _0687_ sky130_fd_sc_hd__a22o_1
X_5382_ _1488_ _1394_ VGND VGND VPWR VPWR 
+ _1582_
+ sky130_fd_sc_hd__or2_1
X_5383_ _1582_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__clkbuf_4
X_5384_ _1583_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__inv_2
X_5385_ \gpio_configure[21][7]\ _1583_ \cdata[7]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0686_ sky130_fd_sc_hd__a22o_1
X_5386_ \gpio_configure[21][6]\ _1583_ \cdata[6]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0685_ sky130_fd_sc_hd__a22o_1
X_5387_ \gpio_configure[21][5]\ _1583_ \cdata[5]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0684_ sky130_fd_sc_hd__a22o_1
X_5388_ \gpio_configure[21][4]\ _1583_ net360 _1584_ VGND VGND 
+ VPWR
+ VPWR _0683_ sky130_fd_sc_hd__a22o_1
X_5389_ \gpio_configure[21][3]\ _1583_ \cdata[3]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0682_ sky130_fd_sc_hd__a22o_1
X_5390_ \gpio_configure[21][2]\ _1583_ \cdata[2]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0681_ sky130_fd_sc_hd__a22o_1
X_5391_ \gpio_configure[21][1]\ _1583_ \cdata[1]\ _1584_ VGND VGND 
+ VPWR
+ VPWR _0680_ sky130_fd_sc_hd__a22o_1
X_5392_ \gpio_configure[21][0]\ _1583_ net368 _1584_ VGND VGND 
+ VPWR
+ VPWR _0679_ sky130_fd_sc_hd__a22o_1
X_5393_ _1488_ _1295_ VGND VGND VPWR VPWR 
+ _1585_
+ sky130_fd_sc_hd__or2_1
X_5394_ _1585_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__clkbuf_4
X_5395_ _1586_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__inv_2
X_5396_ \gpio_configure[31][7]\ _1586_ \cdata[7]\ _1587_ VGND VGND 
+ VPWR
+ VPWR _0678_ sky130_fd_sc_hd__a22o_1
X_5397_ \gpio_configure[31][6]\ _1586_ \cdata[6]\ _1587_ VGND VGND 
+ VPWR
+ VPWR _0677_ sky130_fd_sc_hd__a22o_1
X_5398_ \gpio_configure[31][5]\ _1586_ \cdata[5]\ _1587_ VGND VGND 
+ VPWR
+ VPWR _0676_ sky130_fd_sc_hd__a22o_1
X_5399_ \gpio_configure[31][4]\ _1586_ net359 _1587_ VGND VGND 
+ VPWR
+ VPWR _0675_ sky130_fd_sc_hd__a22o_1
X_5400_ \gpio_configure[31][3]\ _1586_ net361 _1587_ VGND VGND 
+ VPWR
+ VPWR _0674_ sky130_fd_sc_hd__a22o_1
X_5401_ \gpio_configure[31][2]\ _1586_ net363 _1587_ VGND VGND 
+ VPWR
+ VPWR _0673_ sky130_fd_sc_hd__a22o_1
X_5402_ \gpio_configure[31][1]\ _1586_ net366 _1587_ VGND VGND 
+ VPWR
+ VPWR _0672_ sky130_fd_sc_hd__a22o_1
X_5403_ \gpio_configure[31][0]\ _1586_ net368 _1587_ VGND VGND 
+ VPWR
+ VPWR _0671_ sky130_fd_sc_hd__a22o_1
X_5404_ _1551_ _1377_ VGND VGND VPWR VPWR 
+ _1588_
+ sky130_fd_sc_hd__or2_1
X_5405_ _1588_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__clkbuf_2
X_5406_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__inv_2
X_5407_ \gpio_configure[21][12]\ _1589_ net359 _1590_ VGND VGND 
+ VPWR
+ VPWR _0670_ sky130_fd_sc_hd__a22o_1
X_5408_ \gpio_configure[21][11]\ _1589_ net361 _1590_ VGND VGND 
+ VPWR
+ VPWR _0669_ sky130_fd_sc_hd__a22o_1
X_5409_ \gpio_configure[21][10]\ _1589_ net363 _1590_ VGND VGND 
+ VPWR
+ VPWR _0668_ sky130_fd_sc_hd__a22o_1
X_5410_ \gpio_configure[21][9]\ _1589_ net365 _1590_ VGND VGND 
+ VPWR
+ VPWR _0667_ sky130_fd_sc_hd__a22o_1
X_5411_ \gpio_configure[21][8]\ _1589_ net367 _1590_ VGND VGND 
+ VPWR
+ VPWR _0666_ sky130_fd_sc_hd__a22o_1
X_5412_ _1551_ _1380_ VGND VGND VPWR VPWR 
+ _1591_
+ sky130_fd_sc_hd__or2_1
X_5413_ _1591_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__clkbuf_2
X_5414_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__inv_2
X_5415_ \gpio_configure[32][12]\ _1592_ \cdata[4]\ _1593_ VGND VGND 
+ VPWR
+ VPWR _0665_ sky130_fd_sc_hd__a22o_1
X_5416_ \gpio_configure[32][11]\ _1592_ net361 _1593_ VGND VGND 
+ VPWR
+ VPWR _0664_ sky130_fd_sc_hd__a22o_1
X_5417_ \gpio_configure[32][10]\ _1592_ net363 _1593_ VGND VGND 
+ VPWR
+ VPWR _0663_ sky130_fd_sc_hd__a22o_1
X_5418_ \gpio_configure[32][9]\ _1592_ net365 _1593_ VGND VGND 
+ VPWR
+ VPWR _0662_ sky130_fd_sc_hd__a22o_1
X_5419_ \gpio_configure[32][8]\ _1592_ net367 _1593_ VGND VGND 
+ VPWR
+ VPWR _0661_ sky130_fd_sc_hd__a22o_1
X_5420_ _1488_ _1392_ VGND VGND VPWR VPWR 
+ _1594_
+ sky130_fd_sc_hd__or2_1
X_5421_ _1594_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__clkbuf_4
X_5422_ _1595_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__inv_2
X_5423_ \gpio_configure[20][7]\ _1595_ \cdata[7]\ _1596_ VGND VGND 
+ VPWR
+ VPWR _0660_ sky130_fd_sc_hd__a22o_1
X_5424_ \gpio_configure[20][6]\ _1595_ \cdata[6]\ _1596_ VGND VGND 
+ VPWR
+ VPWR _0659_ sky130_fd_sc_hd__a22o_1
X_5425_ \gpio_configure[20][5]\ _1595_ \cdata[5]\ _1596_ VGND VGND 
+ VPWR
+ VPWR _0658_ sky130_fd_sc_hd__a22o_1
X_5426_ \gpio_configure[20][4]\ _1595_ net360 _1596_ VGND VGND 
+ VPWR
+ VPWR _0657_ sky130_fd_sc_hd__a22o_1
X_5427_ \gpio_configure[20][3]\ _1595_ net362 _1596_ VGND VGND 
+ VPWR
+ VPWR _0656_ sky130_fd_sc_hd__a22o_1
X_5428_ \gpio_configure[20][2]\ _1595_ \cdata[2]\ _1596_ VGND VGND 
+ VPWR
+ VPWR _0655_ sky130_fd_sc_hd__a22o_1
X_5429_ \gpio_configure[20][1]\ _1595_ net366 _1596_ VGND VGND 
+ VPWR
+ VPWR _0654_ sky130_fd_sc_hd__a22o_1
X_5430_ \gpio_configure[20][0]\ _1595_ \cdata[0]\ _1596_ VGND VGND 
+ VPWR
+ VPWR _0653_ sky130_fd_sc_hd__a22o_1
X_5431_ _1488_ _1312_ VGND VGND VPWR VPWR 
+ _1597_
+ sky130_fd_sc_hd__or2_1
X_5432_ _1597_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__clkbuf_4
X_5433_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__inv_2
X_5434_ \gpio_configure[32][7]\ _1598_ \cdata[7]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0652_ sky130_fd_sc_hd__a22o_1
X_5435_ \gpio_configure[32][6]\ _1598_ \cdata[6]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0651_ sky130_fd_sc_hd__a22o_1
X_5436_ \gpio_configure[32][5]\ _1598_ \cdata[5]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0650_ sky130_fd_sc_hd__a22o_1
X_5437_ \gpio_configure[32][4]\ _1598_ net360 _1599_ VGND VGND 
+ VPWR
+ VPWR _0649_ sky130_fd_sc_hd__a22o_1
X_5438_ \gpio_configure[32][3]\ _1598_ \cdata[3]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0648_ sky130_fd_sc_hd__a22o_1
X_5439_ \gpio_configure[32][2]\ _1598_ \cdata[2]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0647_ sky130_fd_sc_hd__a22o_1
X_5440_ \gpio_configure[32][1]\ _1598_ \cdata[1]\ _1599_ VGND VGND 
+ VPWR
+ VPWR _0646_ sky130_fd_sc_hd__a22o_1
X_5441_ \gpio_configure[32][0]\ _1598_ net368 _1599_ VGND VGND 
+ VPWR
+ VPWR _0645_ sky130_fd_sc_hd__a22o_1
X_5442_ _1551_ _1327_ VGND VGND VPWR VPWR 
+ _1600_
+ sky130_fd_sc_hd__or2_1
X_5443_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__clkbuf_2
X_5444_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__inv_2
X_5445_ \gpio_configure[20][12]\ _1601_ net359 _1602_ VGND VGND 
+ VPWR
+ VPWR _0644_ sky130_fd_sc_hd__a22o_1
X_5446_ \gpio_configure[20][11]\ _1601_ net361 _1602_ VGND VGND 
+ VPWR
+ VPWR _0643_ sky130_fd_sc_hd__a22o_1
X_5447_ \gpio_configure[20][10]\ _1601_ net363 _1602_ VGND VGND 
+ VPWR
+ VPWR _0642_ sky130_fd_sc_hd__a22o_1
X_5448_ \gpio_configure[20][9]\ _1601_ net365 _1602_ VGND VGND 
+ VPWR
+ VPWR _0641_ sky130_fd_sc_hd__a22o_1
X_5449_ \gpio_configure[20][8]\ _1601_ net367 _1602_ VGND VGND 
+ VPWR
+ VPWR _0640_ sky130_fd_sc_hd__a22o_1
X_5450_ _1551_ _1368_ VGND VGND VPWR VPWR 
+ _1603_
+ sky130_fd_sc_hd__or2_1
X_5451_ _1603_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__buf_2
X_5452_ _1604_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__clkinv_2
X_5453_ \gpio_configure[33][12]\ _1604_ net359 _1605_ VGND VGND 
+ VPWR
+ VPWR _0639_ sky130_fd_sc_hd__a22o_1
X_5454_ \gpio_configure[33][11]\ _1604_ net361 _1605_ VGND VGND 
+ VPWR
+ VPWR _0638_ sky130_fd_sc_hd__a22o_1
X_5455_ \gpio_configure[33][10]\ _1604_ net363 _1605_ VGND VGND 
+ VPWR
+ VPWR _0637_ sky130_fd_sc_hd__a22o_1
X_5456_ \gpio_configure[33][9]\ _1604_ net365 _1605_ VGND VGND 
+ VPWR
+ VPWR _0636_ sky130_fd_sc_hd__a22o_1
X_5457_ \gpio_configure[33][8]\ _1604_ net367 _1605_ VGND VGND 
+ VPWR
+ VPWR _0635_ sky130_fd_sc_hd__a22o_1
X_5458_ _1488_ _1406_ VGND VGND VPWR VPWR 
+ _1606_
+ sky130_fd_sc_hd__or2_1
X_5459_ _1606_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__clkbuf_4
X_5460_ _1607_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__inv_2
X_5461_ \gpio_configure[19][7]\ _1607_ \cdata[7]\ _1608_ VGND VGND 
+ VPWR
+ VPWR _0634_ sky130_fd_sc_hd__a22o_1
X_5462_ \gpio_configure[19][6]\ _1607_ \cdata[6]\ _1608_ VGND VGND 
+ VPWR
+ VPWR _0633_ sky130_fd_sc_hd__a22o_1
X_5463_ \gpio_configure[19][5]\ _1607_ \cdata[5]\ _1608_ VGND VGND 
+ VPWR
+ VPWR _0632_ sky130_fd_sc_hd__a22o_1
X_5464_ \gpio_configure[19][4]\ _1607_ net359 _1608_ VGND VGND 
+ VPWR
+ VPWR _0631_ sky130_fd_sc_hd__a22o_1
X_5465_ \gpio_configure[19][3]\ _1607_ net361 _1608_ VGND VGND 
+ VPWR
+ VPWR _0630_ sky130_fd_sc_hd__a22o_1
X_5466_ \gpio_configure[19][2]\ _1607_ net363 _1608_ VGND VGND 
+ VPWR
+ VPWR _0629_ sky130_fd_sc_hd__a22o_1
X_5467_ \gpio_configure[19][1]\ _1607_ net365 _1608_ VGND VGND 
+ VPWR
+ VPWR _0628_ sky130_fd_sc_hd__a22o_1
X_5468_ \gpio_configure[19][0]\ _1607_ net367 _1608_ VGND VGND 
+ VPWR
+ VPWR _0627_ sky130_fd_sc_hd__a22o_1
X_5469_ _1488_ _1224_ VGND VGND VPWR VPWR 
+ _1609_
+ sky130_fd_sc_hd__or2_1
X_5470_ _1609_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__clkbuf_4
X_5471_ _1610_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__inv_2
X_5472_ \gpio_configure[33][7]\ _1610_ \cdata[7]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0626_ sky130_fd_sc_hd__a22o_1
X_5473_ \gpio_configure[33][6]\ _1610_ \cdata[6]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0625_ sky130_fd_sc_hd__a22o_1
X_5474_ \gpio_configure[33][5]\ _1610_ \cdata[5]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0624_ sky130_fd_sc_hd__a22o_1
X_5475_ \gpio_configure[33][4]\ _1610_ net360 _1611_ VGND VGND 
+ VPWR
+ VPWR _0623_ sky130_fd_sc_hd__a22o_1
X_5476_ \gpio_configure[33][3]\ _1610_ \cdata[3]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0622_ sky130_fd_sc_hd__a22o_1
X_5477_ \gpio_configure[33][2]\ _1610_ \cdata[2]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0621_ sky130_fd_sc_hd__a22o_1
X_5478_ \gpio_configure[33][1]\ _1610_ \cdata[1]\ _1611_ VGND VGND 
+ VPWR
+ VPWR _0620_ sky130_fd_sc_hd__a22o_1
X_5479_ \gpio_configure[33][0]\ _1610_ net368 _1611_ VGND VGND 
+ VPWR
+ VPWR _0619_ sky130_fd_sc_hd__a22o_1
X_5480_ _1551_ _1396_ VGND VGND VPWR VPWR 
+ _1612_
+ sky130_fd_sc_hd__or2_1
X_5481_ _1612_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__clkbuf_2
X_5482_ _1613_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__inv_2
X_5483_ \gpio_configure[19][12]\ _1613_ net359 _1614_ VGND VGND 
+ VPWR
+ VPWR _0618_ sky130_fd_sc_hd__a22o_1
X_5484_ \gpio_configure[19][11]\ _1613_ net361 _1614_ VGND VGND 
+ VPWR
+ VPWR _0617_ sky130_fd_sc_hd__a22o_1
X_5485_ \gpio_configure[19][10]\ _1613_ net363 _1614_ VGND VGND 
+ VPWR
+ VPWR _0616_ sky130_fd_sc_hd__a22o_1
X_5486_ \gpio_configure[19][9]\ _1613_ net365 _1614_ VGND VGND 
+ VPWR
+ VPWR _0615_ sky130_fd_sc_hd__a22o_1
X_5487_ \gpio_configure[19][8]\ _1613_ net367 _1614_ VGND VGND 
+ VPWR
+ VPWR _0614_ sky130_fd_sc_hd__a22o_1
X_5488_ _1551_ _1266_ VGND VGND VPWR VPWR 
+ _1615_
+ sky130_fd_sc_hd__or2_1
X_5489_ _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__clkbuf_2
X_5490_ _1616_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__inv_2
X_5491_ \gpio_configure[34][12]\ _1616_ net359 _1617_ VGND VGND 
+ VPWR
+ VPWR _0613_ sky130_fd_sc_hd__a22o_1
X_5492_ \gpio_configure[34][11]\ _1616_ net361 _1617_ VGND VGND 
+ VPWR
+ VPWR _0612_ sky130_fd_sc_hd__a22o_1
X_5493_ \gpio_configure[34][10]\ _1616_ net363 _1617_ VGND VGND 
+ VPWR
+ VPWR _0611_ sky130_fd_sc_hd__a22o_1
X_5494_ \gpio_configure[34][9]\ _1616_ net365 _1617_ VGND VGND 
+ VPWR
+ VPWR _0610_ sky130_fd_sc_hd__a22o_1
X_5495_ \gpio_configure[34][8]\ _1616_ net367 _1617_ VGND VGND 
+ VPWR
+ VPWR _0609_ sky130_fd_sc_hd__a22o_1
X_5496_ _1488_ _1355_ VGND VGND VPWR VPWR 
+ _1618_
+ sky130_fd_sc_hd__or2_1
X_5497_ _1618_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__clkbuf_4
X_5498_ _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__inv_2
X_5499_ \gpio_configure[18][7]\ _1619_ \cdata[7]\ _1620_ VGND VGND 
+ VPWR
+ VPWR _0608_ sky130_fd_sc_hd__a22o_1
X_5500_ \gpio_configure[18][6]\ _1619_ \cdata[6]\ _1620_ VGND VGND 
+ VPWR
+ VPWR _0607_ sky130_fd_sc_hd__a22o_1
X_5501_ \gpio_configure[18][5]\ _1619_ \cdata[5]\ _1620_ VGND VGND 
+ VPWR
+ VPWR _0606_ sky130_fd_sc_hd__a22o_1
X_5502_ \gpio_configure[18][4]\ _1619_ net360 _1620_ VGND VGND 
+ VPWR
+ VPWR _0605_ sky130_fd_sc_hd__a22o_1
X_5503_ \gpio_configure[18][3]\ _1619_ net362 _1620_ VGND VGND 
+ VPWR
+ VPWR _0604_ sky130_fd_sc_hd__a22o_1
X_5504_ \gpio_configure[18][2]\ _1619_ net364 _1620_ VGND VGND 
+ VPWR
+ VPWR _0603_ sky130_fd_sc_hd__a22o_1
X_5505_ \gpio_configure[18][1]\ _1619_ net366 _1620_ VGND VGND 
+ VPWR
+ VPWR _0602_ sky130_fd_sc_hd__a22o_1
X_5506_ \gpio_configure[18][0]\ _1619_ net368 _1620_ VGND VGND 
+ VPWR
+ VPWR _0601_ sky130_fd_sc_hd__a22o_1
X_5507_ _1488_ _1155_ VGND VGND VPWR VPWR 
+ _1621_
+ sky130_fd_sc_hd__or2_1
X_5508_ _1621_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__clkbuf_4
X_5509_ _1622_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__inv_2
X_5510_ \gpio_configure[34][7]\ _1622_ \cdata[7]\ _1623_ VGND VGND 
+ VPWR
+ VPWR _0600_ sky130_fd_sc_hd__a22o_1
X_5511_ \gpio_configure[34][6]\ _1622_ \cdata[6]\ _1623_ VGND VGND 
+ VPWR
+ VPWR _0599_ sky130_fd_sc_hd__a22o_1
X_5512_ \gpio_configure[34][5]\ _1622_ \cdata[5]\ _1623_ VGND VGND 
+ VPWR
+ VPWR _0598_ sky130_fd_sc_hd__a22o_1
X_5513_ \gpio_configure[34][4]\ _1622_ net360 _1623_ VGND VGND 
+ VPWR
+ VPWR _0597_ sky130_fd_sc_hd__a22o_1
X_5514_ \gpio_configure[34][3]\ _1622_ net362 _1623_ VGND VGND 
+ VPWR
+ VPWR _0596_ sky130_fd_sc_hd__a22o_1
X_5515_ \gpio_configure[34][2]\ _1622_ net364 _1623_ VGND VGND 
+ VPWR
+ VPWR _0595_ sky130_fd_sc_hd__a22o_1
X_5516_ \gpio_configure[34][1]\ _1622_ net366 _1623_ VGND VGND 
+ VPWR
+ VPWR _0594_ sky130_fd_sc_hd__a22o_1
X_5517_ \gpio_configure[34][0]\ _1622_ \cdata[0]\ _1623_ VGND VGND 
+ VPWR
+ VPWR _0593_ sky130_fd_sc_hd__a22o_1
X_5518_ _1551_ _1398_ VGND VGND VPWR VPWR 
+ _1624_
+ sky130_fd_sc_hd__or2_1
X_5519_ _1624_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__clkbuf_2
X_5520_ _1625_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__inv_2
X_5521_ \gpio_configure[18][12]\ _1625_ net359 _1626_ VGND VGND 
+ VPWR
+ VPWR _0592_ sky130_fd_sc_hd__a22o_1
X_5522_ \gpio_configure[18][11]\ _1625_ net361 _1626_ VGND VGND 
+ VPWR
+ VPWR _0591_ sky130_fd_sc_hd__a22o_1
X_5523_ \gpio_configure[18][10]\ _1625_ net363 _1626_ VGND VGND 
+ VPWR
+ VPWR _0590_ sky130_fd_sc_hd__a22o_1
X_5524_ \gpio_configure[18][9]\ _1625_ net365 _1626_ VGND VGND 
+ VPWR
+ VPWR _0589_ sky130_fd_sc_hd__a22o_1
X_5525_ \gpio_configure[18][8]\ _1625_ net367 _1626_ VGND VGND 
+ VPWR
+ VPWR _0588_ sky130_fd_sc_hd__a22o_1
X_5526_ _1551_ _1151_ VGND VGND VPWR VPWR 
+ _1627_
+ sky130_fd_sc_hd__or2_1
X_5527_ _1627_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__clkbuf_2
X_5528_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__inv_2
X_5529_ \gpio_configure[35][12]\ _1628_ \cdata[4]\ _1629_ VGND VGND 
+ VPWR
+ VPWR _0587_ sky130_fd_sc_hd__a22o_1
X_5530_ \gpio_configure[35][11]\ _1628_ \cdata[3]\ _1629_ VGND VGND 
+ VPWR
+ VPWR _0586_ sky130_fd_sc_hd__a22o_1
X_5531_ \gpio_configure[35][10]\ _1628_ \cdata[2]\ _1629_ VGND VGND 
+ VPWR
+ VPWR _0585_ sky130_fd_sc_hd__a22o_1
X_5532_ \gpio_configure[35][9]\ _1628_ net365 _1629_ VGND VGND 
+ VPWR
+ VPWR _0584_ sky130_fd_sc_hd__a22o_1
X_5533_ \gpio_configure[35][8]\ _1628_ \cdata[0]\ _1629_ VGND VGND 
+ VPWR
+ VPWR _0583_ sky130_fd_sc_hd__a22o_1
X_5534_ _1488_ _1284_ VGND VGND VPWR VPWR 
+ _1630_
+ sky130_fd_sc_hd__or2_1
X_5535_ _1630_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__clkbuf_4
X_5536_ _1631_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__inv_2
X_5537_ \gpio_configure[17][7]\ _1631_ \cdata[7]\ _1632_ VGND VGND 
+ VPWR
+ VPWR _0582_ sky130_fd_sc_hd__a22o_1
X_5538_ \gpio_configure[17][6]\ _1631_ \cdata[6]\ _1632_ VGND VGND 
+ VPWR
+ VPWR _0581_ sky130_fd_sc_hd__a22o_1
X_5539_ \gpio_configure[17][5]\ _1631_ \cdata[5]\ _1632_ VGND VGND 
+ VPWR
+ VPWR _0580_ sky130_fd_sc_hd__a22o_1
X_5540_ \gpio_configure[17][4]\ _1631_ net360 _1632_ VGND VGND 
+ VPWR
+ VPWR _0579_ sky130_fd_sc_hd__a22o_1
X_5541_ \gpio_configure[17][3]\ _1631_ net362 _1632_ VGND VGND 
+ VPWR
+ VPWR _0578_ sky130_fd_sc_hd__a22o_1
X_5542_ \gpio_configure[17][2]\ _1631_ net364 _1632_ VGND VGND 
+ VPWR
+ VPWR _0577_ sky130_fd_sc_hd__a22o_1
X_5543_ \gpio_configure[17][1]\ _1631_ net366 _1632_ VGND VGND 
+ VPWR
+ VPWR _0576_ sky130_fd_sc_hd__a22o_1
X_5544_ \gpio_configure[17][0]\ _1631_ net368 _1632_ VGND VGND 
+ VPWR
+ VPWR _0575_ sky130_fd_sc_hd__a22o_1
X_5545_ _1488_ _1231_ VGND VGND VPWR VPWR 
+ _1633_
+ sky130_fd_sc_hd__or2_1
X_5546_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__clkbuf_4
X_5547_ _1634_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__inv_2
X_5548_ \gpio_configure[35][7]\ _1634_ \cdata[7]\ _1635_ VGND VGND 
+ VPWR
+ VPWR _0574_ sky130_fd_sc_hd__a22o_1
X_5549_ \gpio_configure[35][6]\ _1634_ \cdata[6]\ _1635_ VGND VGND 
+ VPWR
+ VPWR _0573_ sky130_fd_sc_hd__a22o_1
X_5550_ \gpio_configure[35][5]\ _1634_ \cdata[5]\ _1635_ VGND VGND 
+ VPWR
+ VPWR _0572_ sky130_fd_sc_hd__a22o_1
X_5551_ \gpio_configure[35][4]\ _1634_ net360 _1635_ VGND VGND 
+ VPWR
+ VPWR _0571_ sky130_fd_sc_hd__a22o_1
X_5552_ \gpio_configure[35][3]\ _1634_ net362 _1635_ VGND VGND 
+ VPWR
+ VPWR _0570_ sky130_fd_sc_hd__a22o_1
X_5553_ \gpio_configure[35][2]\ _1634_ \cdata[2]\ _1635_ VGND VGND 
+ VPWR
+ VPWR _0569_ sky130_fd_sc_hd__a22o_1
X_5554_ \gpio_configure[35][1]\ _1634_ net366 _1635_ VGND VGND 
+ VPWR
+ VPWR _0568_ sky130_fd_sc_hd__a22o_1
X_5555_ \gpio_configure[35][0]\ _1634_ \cdata[0]\ _1635_ VGND VGND 
+ VPWR
+ VPWR _0567_ sky130_fd_sc_hd__a22o_1
X_5556_ _1551_ _1142_ VGND VGND VPWR VPWR 
+ _1636_
+ sky130_fd_sc_hd__or2_1
X_5557_ _1636_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__clkbuf_2
X_5558_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__inv_2
X_5559_ \gpio_configure[17][12]\ _1637_ \cdata[4]\ _1638_ VGND VGND 
+ VPWR
+ VPWR _0566_ sky130_fd_sc_hd__a22o_1
X_5560_ \gpio_configure[17][11]\ _1637_ \cdata[3]\ _1638_ VGND VGND 
+ VPWR
+ VPWR _0565_ sky130_fd_sc_hd__a22o_1
X_5561_ \gpio_configure[17][10]\ _1637_ \cdata[2]\ _1638_ VGND VGND 
+ VPWR
+ VPWR _0564_ sky130_fd_sc_hd__a22o_1
X_5562_ \gpio_configure[17][9]\ _1637_ net366 _1638_ VGND VGND 
+ VPWR
+ VPWR _0563_ sky130_fd_sc_hd__a22o_1
X_5563_ \gpio_configure[17][8]\ _1637_ \cdata[0]\ _1638_ VGND VGND 
+ VPWR
+ VPWR _0562_ sky130_fd_sc_hd__a22o_1
X_5564_ _1551_ _1243_ VGND VGND VPWR VPWR 
+ _1639_
+ sky130_fd_sc_hd__or2_1
X_5565_ _1639_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__clkbuf_2
X_5566_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__inv_2
X_5567_ \gpio_configure[36][12]\ _1640_ net359 _1641_ VGND VGND 
+ VPWR
+ VPWR _0561_ sky130_fd_sc_hd__a22o_1
X_5568_ \gpio_configure[36][11]\ _1640_ net361 _1641_ VGND VGND 
+ VPWR
+ VPWR _0560_ sky130_fd_sc_hd__a22o_1
X_5569_ \gpio_configure[36][10]\ _1640_ net363 _1641_ VGND VGND 
+ VPWR
+ VPWR _0559_ sky130_fd_sc_hd__a22o_1
X_5570_ \gpio_configure[36][9]\ _1640_ net365 _1641_ VGND VGND 
+ VPWR
+ VPWR _0558_ sky130_fd_sc_hd__a22o_1
X_5571_ \gpio_configure[36][8]\ _1640_ net367 _1641_ VGND VGND 
+ VPWR
+ VPWR _0557_ sky130_fd_sc_hd__a22o_1
X_5572_ _1022_ _1222_ VGND VGND VPWR VPWR 
+ _1642_
+ sky130_fd_sc_hd__or2_1
X_5573_ _1642_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__clkbuf_4
X_5574_ _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__inv_2
X_5575_ \gpio_configure[16][7]\ _1643_ \cdata[7]\ _1644_ VGND VGND 
+ VPWR
+ VPWR _0556_ sky130_fd_sc_hd__a22o_1
X_5576_ \gpio_configure[16][6]\ _1643_ \cdata[6]\ _1644_ VGND VGND 
+ VPWR
+ VPWR _0555_ sky130_fd_sc_hd__a22o_1
X_5577_ \gpio_configure[16][5]\ _1643_ \cdata[5]\ _1644_ VGND VGND 
+ VPWR
+ VPWR _0554_ sky130_fd_sc_hd__a22o_1
X_5578_ \gpio_configure[16][4]\ _1643_ net360 _1644_ VGND VGND 
+ VPWR
+ VPWR _0553_ sky130_fd_sc_hd__a22o_1
X_5579_ \gpio_configure[16][3]\ _1643_ net362 _1644_ VGND VGND 
+ VPWR
+ VPWR _0552_ sky130_fd_sc_hd__a22o_1
X_5580_ \gpio_configure[16][2]\ _1643_ net364 _1644_ VGND VGND 
+ VPWR
+ VPWR _0551_ sky130_fd_sc_hd__a22o_1
X_5581_ \gpio_configure[16][1]\ _1643_ net366 _1644_ VGND VGND 
+ VPWR
+ VPWR _0550_ sky130_fd_sc_hd__a22o_1
X_5582_ \gpio_configure[16][0]\ _1643_ net368 _1644_ VGND VGND 
+ VPWR
+ VPWR _0549_ sky130_fd_sc_hd__a22o_1
X_5583_ _1022_ _1251_ VGND VGND VPWR VPWR 
+ _1645_
+ sky130_fd_sc_hd__or2_1
X_5584_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__clkbuf_4
X_5585_ _1646_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__inv_2
X_5586_ \gpio_configure[36][7]\ _1646_ \cdata[7]\ _1647_ VGND VGND 
+ VPWR
+ VPWR _0548_ sky130_fd_sc_hd__a22o_1
X_5587_ \gpio_configure[36][6]\ _1646_ \cdata[6]\ _1647_ VGND VGND 
+ VPWR
+ VPWR _0547_ sky130_fd_sc_hd__a22o_1
X_5588_ \gpio_configure[36][5]\ _1646_ \cdata[5]\ _1647_ VGND VGND 
+ VPWR
+ VPWR _0546_ sky130_fd_sc_hd__a22o_1
X_5589_ \gpio_configure[36][4]\ _1646_ net360 _1647_ VGND VGND 
+ VPWR
+ VPWR _0545_ sky130_fd_sc_hd__a22o_1
X_5590_ \gpio_configure[36][3]\ _1646_ net362 _1647_ VGND VGND 
+ VPWR
+ VPWR _0544_ sky130_fd_sc_hd__a22o_1
X_5591_ \gpio_configure[36][2]\ _1646_ \cdata[2]\ _1647_ VGND VGND 
+ VPWR
+ VPWR _0543_ sky130_fd_sc_hd__a22o_1
X_5592_ \gpio_configure[36][1]\ _1646_ net366 _1647_ VGND VGND 
+ VPWR
+ VPWR _0542_ sky130_fd_sc_hd__a22o_1
X_5593_ \gpio_configure[36][0]\ _1646_ \cdata[0]\ _1647_ VGND VGND 
+ VPWR
+ VPWR _0541_ sky130_fd_sc_hd__a22o_1
X_5594_ _1551_ _1198_ VGND VGND VPWR VPWR 
+ _1648_
+ sky130_fd_sc_hd__or2_1
X_5595_ _1648_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__clkbuf_2
X_5596_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__inv_2
X_5597_ \gpio_configure[16][12]\ _1649_ \cdata[4]\ _1650_ VGND VGND 
+ VPWR
+ VPWR _0540_ sky130_fd_sc_hd__a22o_1
X_5598_ \gpio_configure[16][11]\ _1649_ \cdata[3]\ _1650_ VGND VGND 
+ VPWR
+ VPWR _0539_ sky130_fd_sc_hd__a22o_1
X_5599_ \gpio_configure[16][10]\ _1649_ \cdata[2]\ _1650_ VGND VGND 
+ VPWR
+ VPWR _0538_ sky130_fd_sc_hd__a22o_1
X_5600_ \gpio_configure[16][9]\ _1649_ net366 _1650_ VGND VGND 
+ VPWR
+ VPWR _0537_ sky130_fd_sc_hd__a22o_1
X_5601_ \gpio_configure[16][8]\ _1649_ \cdata[0]\ _1650_ VGND VGND 
+ VPWR
+ VPWR _0536_ sky130_fd_sc_hd__a22o_1
X_5602_ _1551_ _1229_ VGND VGND VPWR VPWR 
+ _1651_
+ sky130_fd_sc_hd__or2_1
X_5603_ _1651_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__clkbuf_2
X_5604_ _1652_ VGND VGND VPWR VPWR _1653_ sky130_fd_sc_hd__inv_2
X_5605_ \gpio_configure[37][12]\ _1652_ \cdata[4]\ _1653_ VGND VGND 
+ VPWR
+ VPWR _0535_ sky130_fd_sc_hd__a22o_1
X_5606_ \gpio_configure[37][11]\ _1652_ net361 _1653_ VGND VGND 
+ VPWR
+ VPWR _0534_ sky130_fd_sc_hd__a22o_1
X_5607_ \gpio_configure[37][10]\ _1652_ net363 _1653_ VGND VGND 
+ VPWR
+ VPWR _0533_ sky130_fd_sc_hd__a22o_1
X_5608_ \gpio_configure[37][9]\ _1652_ net365 _1653_ VGND VGND 
+ VPWR
+ VPWR _0532_ sky130_fd_sc_hd__a22o_1
X_5609_ \gpio_configure[37][8]\ _1652_ net367 _1653_ VGND VGND 
+ VPWR
+ VPWR _0531_ sky130_fd_sc_hd__a22o_1
X_5610_ _1022_ _1239_ VGND VGND VPWR VPWR 
+ _1654_
+ sky130_fd_sc_hd__or2_1
X_5611_ _1654_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__clkbuf_4
X_5612_ _1655_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__clkinv_2
X_5613_ \gpio_configure[15][7]\ _1655_ \cdata[7]\ _1656_ VGND VGND 
+ VPWR
+ VPWR _0530_ sky130_fd_sc_hd__a22o_1
X_5614_ \gpio_configure[15][6]\ _1655_ \cdata[6]\ _1656_ VGND VGND 
+ VPWR
+ VPWR _0529_ sky130_fd_sc_hd__a22o_1
X_5615_ \gpio_configure[15][5]\ _1655_ \cdata[5]\ _1656_ VGND VGND 
+ VPWR
+ VPWR _0528_ sky130_fd_sc_hd__a22o_1
X_5616_ \gpio_configure[15][4]\ _1655_ net360 _1656_ VGND VGND 
+ VPWR
+ VPWR _0527_ sky130_fd_sc_hd__a22o_1
X_5617_ \gpio_configure[15][3]\ _1655_ \cdata[3]\ _1656_ VGND VGND 
+ VPWR
+ VPWR _0526_ sky130_fd_sc_hd__a22o_1
X_5618_ \gpio_configure[15][2]\ _1655_ net364 _1656_ VGND VGND 
+ VPWR
+ VPWR _0525_ sky130_fd_sc_hd__a22o_1
X_5619_ \gpio_configure[15][1]\ _1655_ \cdata[1]\ _1656_ VGND VGND 
+ VPWR
+ VPWR _0524_ sky130_fd_sc_hd__a22o_1
X_5620_ \gpio_configure[15][0]\ _1655_ net368 _1656_ VGND VGND 
+ VPWR
+ VPWR _0523_ sky130_fd_sc_hd__a22o_1
X_5621_ _1022_ _1212_ VGND VGND VPWR VPWR 
+ _1657_
+ sky130_fd_sc_hd__or2_1
X_5622_ _1657_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__clkbuf_4
X_5623_ _1658_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__inv_2
X_5624_ \gpio_configure[37][7]\ _1658_ \cdata[7]\ _1659_ VGND VGND 
+ VPWR
+ VPWR _0522_ sky130_fd_sc_hd__a22o_1
X_5625_ \gpio_configure[37][6]\ _1658_ \cdata[6]\ _1659_ VGND VGND 
+ VPWR
+ VPWR _0521_ sky130_fd_sc_hd__a22o_1
X_5626_ \gpio_configure[37][5]\ _1658_ \cdata[5]\ _1659_ VGND VGND 
+ VPWR
+ VPWR _0520_ sky130_fd_sc_hd__a22o_1
X_5627_ \gpio_configure[37][4]\ _1658_ net360 _1659_ VGND VGND 
+ VPWR
+ VPWR _0519_ sky130_fd_sc_hd__a22o_1
X_5628_ \gpio_configure[37][3]\ _1658_ \cdata[3]\ _1659_ VGND VGND 
+ VPWR
+ VPWR _0518_ sky130_fd_sc_hd__a22o_1
X_5629_ \gpio_configure[37][2]\ _1658_ net364 _1659_ VGND VGND 
+ VPWR
+ VPWR _0517_ sky130_fd_sc_hd__a22o_1
X_5630_ \gpio_configure[37][1]\ _1658_ \cdata[1]\ _1659_ VGND VGND 
+ VPWR
+ VPWR _0516_ sky130_fd_sc_hd__a22o_1
X_5631_ \gpio_configure[37][0]\ _1658_ net368 _1659_ VGND VGND 
+ VPWR
+ VPWR _0515_ sky130_fd_sc_hd__a22o_1
X_5632_ _1551_ _1190_ VGND VGND VPWR VPWR 
+ _1660_
+ sky130_fd_sc_hd__or2_1
X_5633_ _1660_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__clkbuf_2
X_5634_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__inv_2
X_5635_ \gpio_configure[15][12]\ _1661_ \cdata[4]\ _1662_ VGND VGND 
+ VPWR
+ VPWR _0514_ sky130_fd_sc_hd__a22o_1
X_5636_ \gpio_configure[15][11]\ _1661_ \cdata[3]\ _1662_ VGND VGND 
+ VPWR
+ VPWR _0513_ sky130_fd_sc_hd__a22o_1
X_5637_ \gpio_configure[15][10]\ _1661_ \cdata[2]\ _1662_ VGND VGND 
+ VPWR
+ VPWR _0512_ sky130_fd_sc_hd__a22o_1
X_5638_ \gpio_configure[15][9]\ _1661_ \cdata[1]\ _1662_ VGND VGND 
+ VPWR
+ VPWR _0511_ sky130_fd_sc_hd__a22o_1
X_5639_ \gpio_configure[15][8]\ _1661_ \cdata[0]\ _1662_ VGND VGND 
+ VPWR
+ VPWR _0510_ sky130_fd_sc_hd__a22o_1
X_5640_ \xfer_count[2]\ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__inv_2
X_5641_ \xfer_count[0]\ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__inv_2
X_5642_ \xfer_state[1]\ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__inv_2
X_5643_ \xfer_state[3]\ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__inv_2
X_5644_ \xfer_state[2]\ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__clkinv_4
X_5645_ _1665_ _1666_ _1667_ \xfer_state[1]\ net306 VGND 
+ VGND
+ VPWR VPWR _1668_ sky130_fd_sc_hd__a32o_2
X_5646_ \xfer_count[1]\ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__inv_2
X_5647_ _1664_ _1668_ _1669_ VGND VGND VPWR 
+ VPWR
+ _1670_ sky130_fd_sc_hd__or3_2
X_5648_ \xfer_count[3]\ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__inv_2
X_5649_ _1671_ _1663_ \xfer_count[1]\ \xfer_count[0]\ VGND VGND 
+ VPWR
+ VPWR _1672_ sky130_fd_sc_hd__or4_1
X_5650_ \xfer_state[1]\ _1672_ \xfer_state[3]\ VGND VGND VPWR 
+ VPWR
+ _1673_ sky130_fd_sc_hd__a21o_1
X_5651_ _1668_ _1673_ VGND VGND VPWR VPWR 
+ _1674_
+ sky130_fd_sc_hd__or2_2
X_5652_ _1663_ _1670_ _1671_ VGND VGND VPWR 
+ VPWR
+ _1675_ sky130_fd_sc_hd__o21ai_2
X_5653_ _1663_ _1670_ _1671_ _1674_ _1675_ VGND 
+ VGND
+ VPWR VPWR _0509_ sky130_fd_sc_hd__o311a_2
X_5654_ _1663_ _1669_ _1664_ _1673_ VGND VGND 
+ VPWR
+ VPWR _1676_ sky130_fd_sc_hd__o31a_1
X_5655_ _1663_ _1670_ _1668_ _1676_ VGND VGND 
+ VPWR
+ VPWR _0508_ sky130_fd_sc_hd__o2bb2a_2
X_5656_ _1664_ _1668_ _1669_ VGND VGND VPWR 
+ VPWR
+ _1677_ sky130_fd_sc_hd__o21ai_2
X_5657_ \xfer_state[1]\ \xfer_state[3]\ _1667_ _1670_ _1677_ VGND 
+ VGND
+ VPWR VPWR _0507_ sky130_fd_sc_hd__o311a_2
X_5658__14 _1668_ VGND VGND VPWR VPWR net392 sky130_fd_sc_hd__inv_2
X_5659_ _1664_ _1668_ \xfer_count[0]\ net392 _1674_ VGND 
+ VGND
+ VPWR VPWR _0506_ sky130_fd_sc_hd__o221a_2
X_5660_ _1022_ _1206_ VGND VGND VPWR VPWR 
+ _1679_
+ sky130_fd_sc_hd__or2_1
X_5661_ _1679_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__clkbuf_4
X_5662_ _1680_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__inv_2
X_5663_ \gpio_configure[14][7]\ _1680_ \cdata[7]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0505_ sky130_fd_sc_hd__a22o_1
X_5664_ \gpio_configure[14][6]\ _1680_ \cdata[6]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0504_ sky130_fd_sc_hd__a22o_1
X_5665_ \gpio_configure[14][5]\ _1680_ \cdata[5]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0503_ sky130_fd_sc_hd__a22o_1
X_5666_ \gpio_configure[14][4]\ _1680_ net360 _1681_ VGND VGND 
+ VPWR
+ VPWR _0502_ sky130_fd_sc_hd__a22o_1
X_5667_ \gpio_configure[14][3]\ _1680_ net362 _1681_ VGND VGND 
+ VPWR
+ VPWR _0501_ sky130_fd_sc_hd__a22o_1
X_5668_ \gpio_configure[14][2]\ _1680_ \cdata[2]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0500_ sky130_fd_sc_hd__a22o_1
X_5669_ \gpio_configure[14][1]\ _1680_ \cdata[1]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0499_ sky130_fd_sc_hd__a22o_1
X_5670_ \gpio_configure[14][0]\ _1680_ \cdata[0]\ _1681_ VGND VGND 
+ VPWR
+ VPWR _0498_ sky130_fd_sc_hd__a22o_1
X_5671_ _1551_ _1186_ VGND VGND VPWR VPWR 
+ _1682_
+ sky130_fd_sc_hd__or2_1
X_5672_ _1682_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__clkbuf_2
X_5673_ _1683_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__inv_2
X_5674_ \gpio_configure[14][12]\ _1683_ \cdata[4]\ _1684_ VGND VGND 
+ VPWR
+ VPWR _0497_ sky130_fd_sc_hd__a22o_1
X_5675_ \gpio_configure[14][11]\ _1683_ \cdata[3]\ _1684_ VGND VGND 
+ VPWR
+ VPWR _0496_ sky130_fd_sc_hd__a22o_1
X_5676_ \gpio_configure[14][10]\ _1683_ \cdata[2]\ _1684_ VGND VGND 
+ VPWR
+ VPWR _0495_ sky130_fd_sc_hd__a22o_1
X_5677_ \gpio_configure[14][9]\ _1683_ net365 _1684_ VGND VGND 
+ VPWR
+ VPWR _0494_ sky130_fd_sc_hd__a22o_1
X_5678_ \gpio_configure[14][8]\ _1683_ \cdata[0]\ _1684_ VGND VGND 
+ VPWR
+ VPWR _0493_ sky130_fd_sc_hd__a22o_1
X_5679_ _1022_ _1200_ VGND VGND VPWR VPWR 
+ _1685_
+ sky130_fd_sc_hd__or2_1
X_5680_ _1685_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__clkbuf_4
X_5681_ _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__clkinv_2
X_5682_ \gpio_configure[13][7]\ _1686_ \cdata[7]\ _1687_ VGND VGND 
+ VPWR
+ VPWR _0492_ sky130_fd_sc_hd__a22o_1
X_5683_ \gpio_configure[13][6]\ _1686_ \cdata[6]\ _1687_ VGND VGND 
+ VPWR
+ VPWR _0491_ sky130_fd_sc_hd__a22o_1
X_5684_ \gpio_configure[13][5]\ _1686_ \cdata[5]\ _1687_ VGND VGND 
+ VPWR
+ VPWR _0490_ sky130_fd_sc_hd__a22o_1
X_5685_ \gpio_configure[13][4]\ _1686_ net360 _1687_ VGND VGND 
+ VPWR
+ VPWR _0489_ sky130_fd_sc_hd__a22o_1
X_5686_ \gpio_configure[13][3]\ _1686_ \cdata[3]\ _1687_ VGND VGND 
+ VPWR
+ VPWR _0488_ sky130_fd_sc_hd__a22o_1
X_5687_ \gpio_configure[13][2]\ _1686_ net364 _1687_ VGND VGND 
+ VPWR
+ VPWR _0487_ sky130_fd_sc_hd__a22o_1
X_5688_ \gpio_configure[13][1]\ _1686_ \cdata[1]\ _1687_ VGND VGND 
+ VPWR
+ VPWR _0486_ sky130_fd_sc_hd__a22o_1
X_5689_ \gpio_configure[13][0]\ _1686_ net368 _1687_ VGND VGND 
+ VPWR
+ VPWR _0485_ sky130_fd_sc_hd__a22o_1
X_5690_ \xfer_state[0]\ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__inv_2
X_5691_ _1688_ \xfer_state[2]\ VGND VGND VPWR VPWR 
+ _1689_
+ sky130_fd_sc_hd__or2_2
X_5692_ _1689_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__inv_2
X_5693_ \pad_count_1[1]\ \pad_count_1[0]\ VGND VGND VPWR VPWR 
+ _1691_
+ sky130_fd_sc_hd__or2_1
X_5694_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__buf_4
X_5695_ \pad_count_1[3]\ \pad_count_1[2]\ VGND VGND VPWR VPWR 
+ _1693_
+ sky130_fd_sc_hd__or2_4
X_5696_ _1667_ _1692_ _1693_ VGND VGND VPWR 
+ VPWR
+ _1694_ sky130_fd_sc_hd__nor3_1
X_5697_ \pad_count_1[4]\ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__inv_2
X_5698_ _1693_ _1692_ _1695_ VGND VGND VPWR 
+ VPWR
+ _1696_ sky130_fd_sc_hd__or3_1
X_5699_ _1696_ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__buf_8
X_5700_ \pad_count_1[4]\ _1690_ _1694_ _1667_ _1697_ VGND 
+ VGND
+ VPWR VPWR _0484_ sky130_fd_sc_hd__o32a_1
X_5701_ \pad_count_1[2]\ _1692_ _1667_ \pad_count_1[3]\ VGND VGND 
+ VPWR
+ VPWR _1698_ sky130_fd_sc_hd__o31a_1
X_5702_ _1694_ _1698_ _1689_ VGND VGND VPWR 
+ VPWR
+ _0483_ sky130_fd_sc_hd__o21a_1
X_5703_ \pad_count_1[2]\ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__inv_2
X_5704_ _1692_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__inv_2
X_5705_ _1667_ _1692_ _1689_ \pad_count_1[2]\ VGND VGND 
+ VPWR
+ VPWR _1701_ sky130_fd_sc_hd__o211a_1
X_5706_ _1699_ _1700_ \xfer_state[2]\ _1701_ VGND VGND 
+ VPWR
+ VPWR _0482_ sky130_fd_sc_hd__a31o_1
X_5707_ \pad_count_1[1]\ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__inv_2
X_5708_ \pad_count_1[0]\ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__inv_2
X_5709_ _1702_ _1703_ VGND VGND VPWR VPWR 
+ _1704_
+ sky130_fd_sc_hd__or2_4
X_5710_ _1704_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__inv_2
X_5711_ \xfer_state[0]\ \xfer_state[2]\ VGND VGND VPWR VPWR 
+ _1706_
+ sky130_fd_sc_hd__or2_1
X_5712_ _1667_ _1700_ _1705_ \pad_count_1[1]\ _1706_ VGND 
+ VGND
+ VPWR VPWR _0481_ sky130_fd_sc_hd__o32a_1
X_5713_ _1706_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__clkinv_2
X_5714_ _1703_ \xfer_state[2]\ \pad_count_1[0]\ _1707_ VGND VGND 
+ VPWR
+ VPWR _0480_ sky130_fd_sc_hd__a22o_1
X_5715_ \pad_count_2[5]\ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__inv_2
X_5716_ \pad_count_2[4]\ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__inv_2
X_5717_ \pad_count_2[1]\ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__inv_2
X_5718_ \pad_count_2[0]\ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__inv_2
X_5719_ _1710_ _1711_ VGND VGND VPWR VPWR 
+ _1712_
+ sky130_fd_sc_hd__or2_2
X_5720_ \pad_count_2[3]\ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__inv_2
X_5721_ \pad_count_2[2]\ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__inv_2
X_5722_ _1713_ _1714_ VGND VGND VPWR VPWR 
+ _1715_
+ sky130_fd_sc_hd__or2_2
X_5723_ _1712_ _1715_ VGND VGND VPWR VPWR 
+ _1716_
+ sky130_fd_sc_hd__or2_2
X_5724_ _1709_ _1667_ _1716_ VGND VGND VPWR 
+ VPWR
+ _1717_ sky130_fd_sc_hd__nor3_1
X_5725_ \pad_count_2[5]\ _1709_ VGND VGND VPWR VPWR 
+ _1718_
+ sky130_fd_sc_hd__or2_1
X_5726_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__buf_4
X_5727_ _1716_ _1719_ VGND VGND VPWR VPWR 
+ _1720_
+ sky130_fd_sc_hd__or2_1
X_5728_ _1720_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__buf_8
X_5729_ _1708_ _1690_ _1717_ _1667_ _1721_ VGND 
+ VGND
+ VPWR VPWR _1722_ sky130_fd_sc_hd__o32a_1
X_5730_ _1722_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__inv_2
X_5731_ \xfer_state[2]\ _1716_ _1707_ VGND VGND VPWR 
+ VPWR
+ _1723_ sky130_fd_sc_hd__a21oi_1
X_5732_ \pad_count_2[4]\ _1723_ _1717_ VGND VGND VPWR 
+ VPWR
+ _0478_ sky130_fd_sc_hd__o21ba_1
X_5733_ \pad_count_2[3]\ _1714_ _1712_ VGND VGND VPWR 
+ VPWR
+ _1724_ sky130_fd_sc_hd__or3_2
X_5734_ _1713_ _1723_ _1667_ _1724_ VGND VGND 
+ VPWR
+ VPWR _0477_ sky130_fd_sc_hd__o22ai_1
X_5735_ \pad_count_2[1]\ \pad_count_2[0]\ \xfer_state[2]\ \pad_count_2[2]\ VGND VGND 
+ VPWR
+ VPWR _1725_ sky130_fd_sc_hd__a31o_1
X_5736_ _1667_ _1712_ _1714_ _1689_ _1725_ VGND 
+ VGND
+ VPWR VPWR _0476_ sky130_fd_sc_hd__o311a_1
X_5737_ _1710_ \pad_count_2[0]\ VGND VGND VPWR VPWR 
+ _1726_
+ sky130_fd_sc_hd__or2_2
X_5738_ \pad_count_2[1]\ _1711_ VGND VGND VPWR VPWR 
+ _1727_
+ sky130_fd_sc_hd__or2_2
X_5739_ \xfer_state[2]\ _1726_ _1727_ _1710_ _1707_ VGND 
+ VGND
+ VPWR VPWR _1728_ sky130_fd_sc_hd__a32o_1
X_5740_ _1728_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__inv_2
X_5741_ \pad_count_2[0]\ _1706_ _1711_ _1667_ VGND VGND 
+ VPWR
+ VPWR _0474_ sky130_fd_sc_hd__o22a_1
X_5742_ _1023_ _1209_ VGND VGND VPWR VPWR 
+ _1729_
+ sky130_fd_sc_hd__or2_1
X_5743_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__clkbuf_2
X_5744_ _1730_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__inv_2
X_5745_ \gpio_configure[13][12]\ _1730_ \cdata[4]\ _1731_ VGND VGND 
+ VPWR
+ VPWR _0473_ sky130_fd_sc_hd__a22o_1
X_5746_ \gpio_configure[13][11]\ _1730_ \cdata[3]\ _1731_ VGND VGND 
+ VPWR
+ VPWR _0472_ sky130_fd_sc_hd__a22o_1
X_5747_ \gpio_configure[13][10]\ _1730_ \cdata[2]\ _1731_ VGND VGND 
+ VPWR
+ VPWR _0471_ sky130_fd_sc_hd__a22o_1
X_5748_ \gpio_configure[13][9]\ _1730_ net366 _1731_ VGND VGND 
+ VPWR
+ VPWR _0470_ sky130_fd_sc_hd__a22o_1
X_5749_ \gpio_configure[13][8]\ _1730_ \cdata[0]\ _1731_ VGND VGND 
+ VPWR
+ VPWR _0469_ sky130_fd_sc_hd__a22o_1
X_5750_ \xfer_state[3]\ net306 VGND VGND VPWR VPWR 
+ _1732_
+ sky130_fd_sc_hd__nor2_2
X_5751_ \xfer_count[3]\ \xfer_count[2]\ _1669_ \xfer_count[0]\ VGND VGND 
+ VPWR
+ VPWR _1733_ sky130_fd_sc_hd__or4_2
X_5752_ \xfer_count[3]\ \xfer_count[2]\ \xfer_count[1]\ VGND VGND VPWR 
+ VPWR
+ _1734_ sky130_fd_sc_hd__or3_1
X_5753_ \xfer_state[3]\ _1733_ _1734_ VGND VGND VPWR 
+ VPWR
+ _1735_ sky130_fd_sc_hd__and3_1
X_5754_ _1665_ _1666_ _1707_ _1735_ VGND VGND 
+ VPWR
+ VPWR _1736_ sky130_fd_sc_hd__a31o_1
X_5755_ _1736_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__inv_2
X_5756_ _1707_ _1732_ _1737_ serial_clock_pre _1736_ VGND 
+ VGND
+ VPWR VPWR _0468_ sky130_fd_sc_hd__a32o_2
X_5757_ _1022_ _1259_ VGND VGND VPWR VPWR 
+ _1738_
+ sky130_fd_sc_hd__or2_1
X_5758_ _1738_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__clkbuf_4
X_5759_ _1739_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__inv_2
X_5760_ \gpio_configure[12][7]\ _1739_ \cdata[7]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0467_ sky130_fd_sc_hd__a22o_1
X_5761_ \gpio_configure[12][6]\ _1739_ \cdata[6]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0466_ sky130_fd_sc_hd__a22o_1
X_5762_ \gpio_configure[12][5]\ _1739_ \cdata[5]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0465_ sky130_fd_sc_hd__a22o_1
X_5763_ \gpio_configure[12][4]\ _1739_ net360 _1740_ VGND VGND 
+ VPWR
+ VPWR _0464_ sky130_fd_sc_hd__a22o_1
X_5764_ \gpio_configure[12][3]\ _1739_ net362 _1740_ VGND VGND 
+ VPWR
+ VPWR _0463_ sky130_fd_sc_hd__a22o_1
X_5765_ \gpio_configure[12][2]\ _1739_ \cdata[2]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0462_ sky130_fd_sc_hd__a22o_1
X_5766_ \gpio_configure[12][1]\ _1739_ \cdata[1]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0461_ sky130_fd_sc_hd__a22o_1
X_5767_ \gpio_configure[12][0]\ _1739_ \cdata[0]\ _1740_ VGND VGND 
+ VPWR
+ VPWR _0460_ sky130_fd_sc_hd__a22o_1
X_5768_ _1023_ _1202_ VGND VGND VPWR VPWR 
+ _1741_
+ sky130_fd_sc_hd__or2_1
X_5769_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__clkbuf_2
X_5770_ _1742_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__inv_2
X_5771_ \gpio_configure[12][12]\ _1742_ net359 _1743_ VGND VGND 
+ VPWR
+ VPWR _0459_ sky130_fd_sc_hd__a22o_1
X_5772_ \gpio_configure[12][11]\ _1742_ net361 _1743_ VGND VGND 
+ VPWR
+ VPWR _0458_ sky130_fd_sc_hd__a22o_1
X_5773_ \gpio_configure[12][10]\ _1742_ net363 _1743_ VGND VGND 
+ VPWR
+ VPWR _0457_ sky130_fd_sc_hd__a22o_1
X_5774_ \gpio_configure[12][9]\ _1742_ net365 _1743_ VGND VGND 
+ VPWR
+ VPWR _0456_ sky130_fd_sc_hd__a22o_1
X_5775_ \gpio_configure[12][8]\ _1742_ net367 _1743_ VGND VGND 
+ VPWR
+ VPWR _0455_ sky130_fd_sc_hd__a22o_1
X_5776_ _1022_ _1188_ VGND VGND VPWR VPWR 
+ _1744_
+ sky130_fd_sc_hd__or2_1
X_5777_ _1744_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__clkbuf_4
X_5778_ _1745_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__clkinv_2
X_5779_ \gpio_configure[11][7]\ _1745_ \cdata[7]\ _1746_ VGND VGND 
+ VPWR
+ VPWR _0454_ sky130_fd_sc_hd__a22o_1
X_5780_ \gpio_configure[11][6]\ _1745_ \cdata[6]\ _1746_ VGND VGND 
+ VPWR
+ VPWR _0453_ sky130_fd_sc_hd__a22o_1
X_5781_ \gpio_configure[11][5]\ _1745_ \cdata[5]\ _1746_ VGND VGND 
+ VPWR
+ VPWR _0452_ sky130_fd_sc_hd__a22o_1
X_5782_ \gpio_configure[11][4]\ _1745_ net360 _1746_ VGND VGND 
+ VPWR
+ VPWR _0451_ sky130_fd_sc_hd__a22o_1
X_5783_ \gpio_configure[11][3]\ _1745_ net362 _1746_ VGND VGND 
+ VPWR
+ VPWR _0450_ sky130_fd_sc_hd__a22o_1
X_5784_ \gpio_configure[11][2]\ _1745_ net364 _1746_ VGND VGND 
+ VPWR
+ VPWR _0449_ sky130_fd_sc_hd__a22o_1
X_5785_ \gpio_configure[11][1]\ _1745_ net366 _1746_ VGND VGND 
+ VPWR
+ VPWR _0448_ sky130_fd_sc_hd__a22o_1
X_5786_ \gpio_configure[11][0]\ _1745_ net368 _1746_ VGND VGND 
+ VPWR
+ VPWR _0447_ sky130_fd_sc_hd__a22o_1
X_5787_ _1734_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__inv_2
X_5788_ \xfer_count[0]\ \xfer_state[3]\ _1747_ serial_load_pre _1736_ VGND 
+ VGND
+ VPWR VPWR _0446_ sky130_fd_sc_hd__a32o_1
X_5789_ _1023_ _1192_ VGND VGND VPWR VPWR 
+ _1748_
+ sky130_fd_sc_hd__or2_1
X_5790_ _1748_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__clkbuf_2
X_5791_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__inv_2
X_5792_ \gpio_configure[11][12]\ _1749_ net359 _1750_ VGND VGND 
+ VPWR
+ VPWR _0445_ sky130_fd_sc_hd__a22o_1
X_5793_ \gpio_configure[11][11]\ _1749_ net361 _1750_ VGND VGND 
+ VPWR
+ VPWR _0444_ sky130_fd_sc_hd__a22o_1
X_5794_ \gpio_configure[11][10]\ _1749_ net363 _1750_ VGND VGND 
+ VPWR
+ VPWR _0443_ sky130_fd_sc_hd__a22o_1
X_5795_ \gpio_configure[11][9]\ _1749_ net366 _1750_ VGND VGND 
+ VPWR
+ VPWR _0442_ sky130_fd_sc_hd__a22o_1
X_5796_ \gpio_configure[11][8]\ _1749_ net367 _1750_ VGND VGND 
+ VPWR
+ VPWR _0441_ sky130_fd_sc_hd__a22o_1
X_5797_ _1022_ _1214_ VGND VGND VPWR VPWR 
+ _1751_
+ sky130_fd_sc_hd__or2_1
X_5798_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__clkbuf_4
X_5799_ _1752_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__clkinv_2
X_5800_ \gpio_configure[10][7]\ _1752_ \cdata[7]\ _1753_ VGND VGND 
+ VPWR
+ VPWR _0440_ sky130_fd_sc_hd__a22o_1
X_5801_ \gpio_configure[10][6]\ _1752_ \cdata[6]\ _1753_ VGND VGND 
+ VPWR
+ VPWR _0439_ sky130_fd_sc_hd__a22o_1
X_5802_ \gpio_configure[10][5]\ _1752_ \cdata[5]\ _1753_ VGND VGND 
+ VPWR
+ VPWR _0438_ sky130_fd_sc_hd__a22o_1
X_5803_ \gpio_configure[10][4]\ _1752_ net360 _1753_ VGND VGND 
+ VPWR
+ VPWR _0437_ sky130_fd_sc_hd__a22o_1
X_5804_ \gpio_configure[10][3]\ _1752_ \cdata[3]\ _1753_ VGND VGND 
+ VPWR
+ VPWR _0436_ sky130_fd_sc_hd__a22o_1
X_5805_ \gpio_configure[10][2]\ _1752_ net364 _1753_ VGND VGND 
+ VPWR
+ VPWR _0435_ sky130_fd_sc_hd__a22o_1
X_5806_ \gpio_configure[10][1]\ _1752_ net366 _1753_ VGND VGND 
+ VPWR
+ VPWR _0434_ sky130_fd_sc_hd__a22o_1
X_5807_ \gpio_configure[10][0]\ _1752_ net368 _1753_ VGND VGND 
+ VPWR
+ VPWR _0433_ sky130_fd_sc_hd__a22o_1
X_5808_ \xfer_state[3]\ _1688_ _1666_ _1733_ serial_busy VGND 
+ VGND
+ VPWR VPWR _1754_ sky130_fd_sc_hd__o221a_1
X_5809_ \xfer_state[0]\ serial_xfer _1666_ _1754_ VGND VGND 
+ VPWR
+ VPWR _0432_ sky130_fd_sc_hd__a31o_1
X_5810_ _1023_ _1165_ VGND VGND VPWR VPWR 
+ _1755_
+ sky130_fd_sc_hd__or2_1
X_5811_ _1755_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__clkbuf_2
X_5812_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__inv_2
X_5813_ \gpio_configure[10][12]\ _1756_ \cdata[4]\ _1757_ VGND VGND 
+ VPWR
+ VPWR _0431_ sky130_fd_sc_hd__a22o_1
X_5814_ \gpio_configure[10][11]\ _1756_ net361 _1757_ VGND VGND 
+ VPWR
+ VPWR _0430_ sky130_fd_sc_hd__a22o_1
X_5815_ \gpio_configure[10][10]\ _1756_ \cdata[2]\ _1757_ VGND VGND 
+ VPWR
+ VPWR _0429_ sky130_fd_sc_hd__a22o_1
X_5816_ \gpio_configure[10][9]\ _1756_ net365 _1757_ VGND VGND 
+ VPWR
+ VPWR _0428_ sky130_fd_sc_hd__a22o_1
X_5817_ \gpio_configure[10][8]\ _1756_ \cdata[0]\ _1757_ VGND VGND 
+ VPWR
+ VPWR _0427_ sky130_fd_sc_hd__a22o_1
X_5818_ _1022_ _1220_ VGND VGND VPWR VPWR 
+ _1758_
+ sky130_fd_sc_hd__or2_1
X_5819_ _1758_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__clkbuf_4
X_5820_ _1759_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__inv_2
X_5821_ \gpio_configure[9][7]\ _1759_ \cdata[7]\ _1760_ VGND VGND 
+ VPWR
+ VPWR _0426_ sky130_fd_sc_hd__a22o_1
X_5822_ \gpio_configure[9][6]\ _1759_ \cdata[6]\ _1760_ VGND VGND 
+ VPWR
+ VPWR _0425_ sky130_fd_sc_hd__a22o_1
X_5823_ \gpio_configure[9][5]\ _1759_ \cdata[5]\ _1760_ VGND VGND 
+ VPWR
+ VPWR _0424_ sky130_fd_sc_hd__a22o_1
X_5824_ \gpio_configure[9][4]\ _1759_ net360 _1760_ VGND VGND 
+ VPWR
+ VPWR _0423_ sky130_fd_sc_hd__a22o_1
X_5825_ \gpio_configure[9][3]\ _1759_ net362 _1760_ VGND VGND 
+ VPWR
+ VPWR _0422_ sky130_fd_sc_hd__a22o_1
X_5826_ \gpio_configure[9][2]\ _1759_ net364 _1760_ VGND VGND 
+ VPWR
+ VPWR _0421_ sky130_fd_sc_hd__a22o_1
X_5827_ \gpio_configure[9][1]\ _1759_ net366 _1760_ VGND VGND 
+ VPWR
+ VPWR _0420_ sky130_fd_sc_hd__a22o_1
X_5828_ \gpio_configure[9][0]\ _1759_ net368 _1760_ VGND VGND 
+ VPWR
+ VPWR _0419_ sky130_fd_sc_hd__a22o_1
X_5829_ _1023_ _1241_ VGND VGND VPWR VPWR 
+ _1761_
+ sky130_fd_sc_hd__or2_1
X_5830_ _1761_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__clkbuf_2
X_5831_ _1762_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__inv_2
X_5832_ \gpio_configure[9][12]\ _1762_ net359 _1763_ VGND VGND 
+ VPWR
+ VPWR _0418_ sky130_fd_sc_hd__a22o_1
X_5833_ \gpio_configure[9][11]\ _1762_ net361 _1763_ VGND VGND 
+ VPWR
+ VPWR _0417_ sky130_fd_sc_hd__a22o_1
X_5834_ \gpio_configure[9][10]\ _1762_ net363 _1763_ VGND VGND 
+ VPWR
+ VPWR _0416_ sky130_fd_sc_hd__a22o_1
X_5835_ \gpio_configure[9][9]\ _1762_ net365 _1763_ VGND VGND 
+ VPWR
+ VPWR _0415_ sky130_fd_sc_hd__a22o_1
X_5836_ \gpio_configure[9][8]\ _1762_ net367 _1763_ VGND VGND 
+ VPWR
+ VPWR _0414_ sky130_fd_sc_hd__a22o_1
X_5837_ _1022_ _1196_ VGND VGND VPWR VPWR 
+ _1764_
+ sky130_fd_sc_hd__or2_1
X_5838_ _1764_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__clkbuf_4
X_5839_ _1765_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__inv_2
X_5840_ \gpio_configure[8][7]\ _1765_ \cdata[7]\ _1766_ VGND VGND 
+ VPWR
+ VPWR _0413_ sky130_fd_sc_hd__a22o_1
X_5841_ \gpio_configure[8][6]\ _1765_ \cdata[6]\ _1766_ VGND VGND 
+ VPWR
+ VPWR _0412_ sky130_fd_sc_hd__a22o_1
X_5842_ \gpio_configure[8][5]\ _1765_ \cdata[5]\ _1766_ VGND VGND 
+ VPWR
+ VPWR _0411_ sky130_fd_sc_hd__a22o_1
X_5843_ \gpio_configure[8][4]\ _1765_ net360 _1766_ VGND VGND 
+ VPWR
+ VPWR _0410_ sky130_fd_sc_hd__a22o_1
X_5844_ \gpio_configure[8][3]\ _1765_ net362 _1766_ VGND VGND 
+ VPWR
+ VPWR _0409_ sky130_fd_sc_hd__a22o_1
X_5845_ \gpio_configure[8][2]\ _1765_ net364 _1766_ VGND VGND 
+ VPWR
+ VPWR _0408_ sky130_fd_sc_hd__a22o_1
X_5846_ \gpio_configure[8][1]\ _1765_ net366 _1766_ VGND VGND 
+ VPWR
+ VPWR _0407_ sky130_fd_sc_hd__a22o_1
X_5847_ \gpio_configure[8][0]\ _1765_ net368 _1766_ VGND VGND 
+ VPWR
+ VPWR _0406_ sky130_fd_sc_hd__a22o_1
X_5848__10 _0042_ VGND VGND VPWR VPWR net388 sky130_fd_sc_hd__inv_4
X_5848__11 _0042_ VGND VGND VPWR VPWR net389 sky130_fd_sc_hd__inv_4
X_5848__12 _0042_ VGND VGND VPWR VPWR net390 sky130_fd_sc_hd__inv_4
X_5848__4 _0042_ VGND VGND VPWR VPWR net382 sky130_fd_sc_hd__inv_4
X_5848__5 _0042_ VGND VGND VPWR VPWR net383 sky130_fd_sc_hd__inv_4
X_5848__6 _0042_ VGND VGND VPWR VPWR net384 sky130_fd_sc_hd__inv_4
X_5848__7 _0042_ VGND VGND VPWR VPWR net385 sky130_fd_sc_hd__inv_4
X_5848__8 _0042_ VGND VGND VPWR VPWR net386 sky130_fd_sc_hd__inv_4
X_5848__9 _0042_ VGND VGND VPWR VPWR net387 sky130_fd_sc_hd__inv_4
X_5849_ net390 VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__buf_1
X_5850_ \serial_data_staging_1[12]\ _0042_ _0002_ _1768_ VGND VGND 
+ VPWR
+ VPWR _0405_ sky130_fd_sc_hd__o22a_2
X_5851_ _1768_ _0001_ _0042_ \serial_data_staging_1[11]\ VGND VGND 
+ VPWR
+ VPWR _0404_ sky130_fd_sc_hd__o22a_2
X_5852_ _1768_ _0000_ _0042_ \serial_data_staging_1[10]\ VGND VGND 
+ VPWR
+ VPWR _0403_ sky130_fd_sc_hd__o22a_2
X_5853_ _1768_ _0011_ _0042_ \serial_data_staging_1[9]\ VGND VGND 
+ VPWR
+ VPWR _0402_ sky130_fd_sc_hd__o22a_2
X_5854_ _1768_ _0010_ _0042_ \serial_data_staging_1[8]\ VGND VGND 
+ VPWR
+ VPWR _0401_ sky130_fd_sc_hd__o22a_2
X_5855_ _1768_ _0009_ _0042_ \serial_data_staging_1[7]\ VGND VGND 
+ VPWR
+ VPWR _0400_ sky130_fd_sc_hd__o22a_2
X_5856_ _1768_ _0008_ _0042_ \serial_data_staging_1[6]\ VGND VGND 
+ VPWR
+ VPWR _0399_ sky130_fd_sc_hd__o22a_2
X_5857_ _1768_ _0007_ _0042_ \serial_data_staging_1[5]\ VGND VGND 
+ VPWR
+ VPWR _0398_ sky130_fd_sc_hd__o22a_2
X_5858_ _1768_ _0006_ _0042_ \serial_data_staging_1[4]\ VGND VGND 
+ VPWR
+ VPWR _0397_ sky130_fd_sc_hd__o22a_2
X_5859_ _1768_ _0005_ _0042_ \serial_data_staging_1[3]\ VGND VGND 
+ VPWR
+ VPWR _0396_ sky130_fd_sc_hd__o22a_2
X_5860_ _1768_ _0004_ _0042_ \serial_data_staging_1[2]\ VGND VGND 
+ VPWR
+ VPWR _0395_ sky130_fd_sc_hd__o22a_2
X_5861_ _1768_ _0003_ _0042_ \serial_data_staging_1[1]\ VGND VGND 
+ VPWR
+ VPWR _0394_ sky130_fd_sc_hd__o22a_2
X_5862_ _0129_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__inv_2
X_5863_ _0042_ _1665_ _1769_ net389 \serial_data_staging_1[0]\ VGND 
+ VGND
+ VPWR VPWR _0393_ sky130_fd_sc_hd__a32o_2
X_5864_ _1023_ _1174_ VGND VGND VPWR VPWR 
+ _1770_
+ sky130_fd_sc_hd__or2_1
X_5865_ _1770_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__clkbuf_2
X_5866_ _1771_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__inv_2
X_5867_ \gpio_configure[8][12]\ _1771_ \cdata[4]\ _1772_ VGND VGND 
+ VPWR
+ VPWR _0392_ sky130_fd_sc_hd__a22o_1
X_5868_ \gpio_configure[8][11]\ _1771_ \cdata[3]\ _1772_ VGND VGND 
+ VPWR
+ VPWR _0391_ sky130_fd_sc_hd__a22o_1
X_5869_ \gpio_configure[8][10]\ _1771_ \cdata[2]\ _1772_ VGND VGND 
+ VPWR
+ VPWR _0390_ sky130_fd_sc_hd__a22o_1
X_5870_ \gpio_configure[8][9]\ _1771_ net365 _1772_ VGND VGND 
+ VPWR
+ VPWR _0389_ sky130_fd_sc_hd__a22o_1
X_5871_ \gpio_configure[8][8]\ _1771_ \cdata[0]\ _1772_ VGND VGND 
+ VPWR
+ VPWR _0388_ sky130_fd_sc_hd__a22o_1
X_5872_ _1022_ _1149_ VGND VGND VPWR VPWR 
+ _1773_
+ sky130_fd_sc_hd__or2_1
X_5873_ _1773_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__clkbuf_4
X_5874_ _1774_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__inv_2
X_5875_ \gpio_configure[7][7]\ _1774_ \cdata[7]\ _1775_ VGND VGND 
+ VPWR
+ VPWR _0387_ sky130_fd_sc_hd__a22o_1
X_5876_ \gpio_configure[7][6]\ _1774_ \cdata[6]\ _1775_ VGND VGND 
+ VPWR
+ VPWR _0386_ sky130_fd_sc_hd__a22o_1
X_5877_ \gpio_configure[7][5]\ _1774_ \cdata[5]\ _1775_ VGND VGND 
+ VPWR
+ VPWR _0385_ sky130_fd_sc_hd__a22o_1
X_5878_ \gpio_configure[7][4]\ _1774_ net360 _1775_ VGND VGND 
+ VPWR
+ VPWR _0384_ sky130_fd_sc_hd__a22o_1
X_5879_ \gpio_configure[7][3]\ _1774_ net362 _1775_ VGND VGND 
+ VPWR
+ VPWR _0383_ sky130_fd_sc_hd__a22o_1
X_5880_ \gpio_configure[7][2]\ _1774_ net364 _1775_ VGND VGND 
+ VPWR
+ VPWR _0382_ sky130_fd_sc_hd__a22o_1
X_5881_ \gpio_configure[7][1]\ _1774_ net366 _1775_ VGND VGND 
+ VPWR
+ VPWR _0381_ sky130_fd_sc_hd__a22o_1
X_5882_ \gpio_configure[7][0]\ _1774_ net368 _1775_ VGND VGND 
+ VPWR
+ VPWR _0380_ sky130_fd_sc_hd__a22o_1
X_5883_ _1768_ _0014_ _0042_ \serial_data_staging_2[12]\ VGND VGND 
+ VPWR
+ VPWR _0379_ sky130_fd_sc_hd__o22a_2
X_5884_ _1768_ _0013_ _0042_ \serial_data_staging_2[11]\ VGND VGND 
+ VPWR
+ VPWR _0378_ sky130_fd_sc_hd__o22a_2
X_5885_ _1768_ _0012_ _0042_ \serial_data_staging_2[10]\ VGND VGND 
+ VPWR
+ VPWR _0377_ sky130_fd_sc_hd__o22a_2
X_5886_ _1768_ _0023_ _0042_ \serial_data_staging_2[9]\ VGND VGND 
+ VPWR
+ VPWR _0376_ sky130_fd_sc_hd__o22a_2
X_5887_ _1768_ _0022_ _0042_ \serial_data_staging_2[8]\ VGND VGND 
+ VPWR
+ VPWR _0375_ sky130_fd_sc_hd__o22a_2
X_5888_ _1768_ _0021_ _0042_ \serial_data_staging_2[7]\ VGND VGND 
+ VPWR
+ VPWR _0374_ sky130_fd_sc_hd__o22a_2
X_5889_ net388 _0020_ _0042_ \serial_data_staging_2[6]\ VGND VGND 
+ VPWR
+ VPWR _0373_ sky130_fd_sc_hd__o22a_2
X_5890_ net387 _0019_ _0042_ \serial_data_staging_2[5]\ VGND VGND 
+ VPWR
+ VPWR _0372_ sky130_fd_sc_hd__o22a_2
X_5891_ net386 _0018_ _0042_ \serial_data_staging_2[4]\ VGND VGND 
+ VPWR
+ VPWR _0371_ sky130_fd_sc_hd__o22a_2
X_5892_ net385 _0017_ _0042_ \serial_data_staging_2[3]\ VGND VGND 
+ VPWR
+ VPWR _0370_ sky130_fd_sc_hd__o22a_2
X_5893_ net384 _0016_ _0042_ \serial_data_staging_2[2]\ VGND VGND 
+ VPWR
+ VPWR _0369_ sky130_fd_sc_hd__o22a_2
X_5894_ net383 _0015_ _0042_ \serial_data_staging_2[1]\ VGND VGND 
+ VPWR
+ VPWR _0368_ sky130_fd_sc_hd__o22a_2
X_5895_ _0102_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__inv_2
X_5896_ _0042_ _1665_ _1776_ net382 \serial_data_staging_2[0]\ VGND 
+ VGND
+ VPWR VPWR _0367_ sky130_fd_sc_hd__a32o_2
X_5897_ _1023_ _1179_ VGND VGND VPWR VPWR 
+ _1777_
+ sky130_fd_sc_hd__or2_1
X_5898_ _1777_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__clkbuf_2
X_5899_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__inv_2
X_5900_ \gpio_configure[7][12]\ _1778_ \cdata[4]\ _1779_ VGND VGND 
+ VPWR
+ VPWR _0366_ sky130_fd_sc_hd__a22o_1
X_5901_ \gpio_configure[7][11]\ _1778_ \cdata[3]\ _1779_ VGND VGND 
+ VPWR
+ VPWR _0365_ sky130_fd_sc_hd__a22o_1
X_5902_ \gpio_configure[7][10]\ _1778_ \cdata[2]\ _1779_ VGND VGND 
+ VPWR
+ VPWR _0364_ sky130_fd_sc_hd__a22o_1
X_5903_ \gpio_configure[7][9]\ _1778_ net365 _1779_ VGND VGND 
+ VPWR
+ VPWR _0363_ sky130_fd_sc_hd__a22o_1
X_5904_ \gpio_configure[7][8]\ _1778_ \cdata[0]\ _1779_ VGND VGND 
+ VPWR
+ VPWR _0362_ sky130_fd_sc_hd__a22o_1
X_5905_ _1022_ _1146_ VGND VGND VPWR VPWR 
+ _1780_
+ sky130_fd_sc_hd__or2_1
X_5906_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__clkbuf_4
X_5907_ _1781_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__inv_2
X_5908_ \gpio_configure[6][7]\ _1781_ \cdata[7]\ _1782_ VGND VGND 
+ VPWR
+ VPWR _0361_ sky130_fd_sc_hd__a22o_1
X_5909_ \gpio_configure[6][6]\ _1781_ \cdata[6]\ _1782_ VGND VGND 
+ VPWR
+ VPWR _0360_ sky130_fd_sc_hd__a22o_1
X_5910_ \gpio_configure[6][5]\ _1781_ \cdata[5]\ _1782_ VGND VGND 
+ VPWR
+ VPWR _0359_ sky130_fd_sc_hd__a22o_1
X_5911_ \gpio_configure[6][4]\ _1781_ net360 _1782_ VGND VGND 
+ VPWR
+ VPWR _0358_ sky130_fd_sc_hd__a22o_1
X_5912_ \gpio_configure[6][3]\ _1781_ net362 _1782_ VGND VGND 
+ VPWR
+ VPWR _0357_ sky130_fd_sc_hd__a22o_1
X_5913_ \gpio_configure[6][2]\ _1781_ net364 _1782_ VGND VGND 
+ VPWR
+ VPWR _0356_ sky130_fd_sc_hd__a22o_1
X_5914_ \gpio_configure[6][1]\ _1781_ net366 _1782_ VGND VGND 
+ VPWR
+ VPWR _0355_ sky130_fd_sc_hd__a22o_1
X_5915_ \gpio_configure[6][0]\ _1781_ net368 _1782_ VGND VGND 
+ VPWR
+ VPWR _0354_ sky130_fd_sc_hd__a22o_1
X_5916_ _1023_ _1255_ VGND VGND VPWR VPWR 
+ _1783_
+ sky130_fd_sc_hd__or2_1
X_5917_ _1783_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__clkbuf_2
X_5918_ _1784_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__inv_2
X_5919_ \gpio_configure[6][12]\ _1784_ net359 _1785_ VGND VGND 
+ VPWR
+ VPWR _0353_ sky130_fd_sc_hd__a22o_1
X_5920_ \gpio_configure[6][11]\ _1784_ net361 _1785_ VGND VGND 
+ VPWR
+ VPWR _0352_ sky130_fd_sc_hd__a22o_1
X_5921_ \gpio_configure[6][10]\ _1784_ net363 _1785_ VGND VGND 
+ VPWR
+ VPWR _0351_ sky130_fd_sc_hd__a22o_1
X_5922_ \gpio_configure[6][9]\ _1784_ net366 _1785_ VGND VGND 
+ VPWR
+ VPWR _0350_ sky130_fd_sc_hd__a22o_1
X_5923_ \gpio_configure[6][8]\ _1784_ net367 _1785_ VGND VGND 
+ VPWR
+ VPWR _0349_ sky130_fd_sc_hd__a22o_1
X_5924_ \wbbd_state[1]\ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__inv_2
X_5925_ net141 net140 net147 net148 VGND VGND 
+ VPWR
+ VPWR _1787_ sky130_fd_sc_hd__or4b_1
X_5926_ net137 net136 net139 net138 VGND VGND 
+ VPWR
+ VPWR _1788_ sky130_fd_sc_hd__or4_1
X_5927_ net133 net132 net135 net134 VGND VGND 
+ VPWR
+ VPWR _1789_ sky130_fd_sc_hd__or4_1
X_5928_ net162 net161 _1789_ VGND VGND VPWR 
+ VPWR
+ _1790_ sky130_fd_sc_hd__or3_1
X_5929_ net146 net145 VGND VGND VPWR VPWR 
+ _1791_
+ sky130_fd_sc_hd__or2_1
X_5930_ net150 net151 net149 net152 VGND VGND 
+ VPWR
+ VPWR _1792_ sky130_fd_sc_hd__or4bb_1
X_5931_ net155 net154 net163 net201 VGND VGND 
+ VPWR
+ VPWR _1793_ sky130_fd_sc_hd__or4bb_1
X_5932_ net144 VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__inv_2
X_5933_ net143 VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__inv_2
X_5934_ _1794_ _1795_ VGND VGND VPWR VPWR 
+ _1796_
+ sky130_fd_sc_hd__or2_1
X_5935_ _1791_ _1792_ _1793_ _1796_ VGND VGND 
+ VPWR
+ VPWR _1797_ sky130_fd_sc_hd__or4b_1
X_5936_ _1787_ _1788_ _1790_ _1797_ VGND VGND 
+ VPWR
+ VPWR _1798_ sky130_fd_sc_hd__or4_2
X_5937_ \wbbd_state[0]\ _1798_ VGND VGND VPWR VPWR 
+ _1799_
+ sky130_fd_sc_hd__and2_1
X_5938_ _1786_ _1799_ VGND VGND VPWR VPWR 
+ _1800_
+ sky130_fd_sc_hd__nor2_1
X_5939_ _1519_ _1798_ VGND VGND VPWR VPWR 
+ _1801_
+ sky130_fd_sc_hd__or2_1
X_5940_ \wbbd_state[0]\ _1080_ net326 _1800_ _1801_ VGND 
+ VGND
+ VPWR VPWR _0348_ sky130_fd_sc_hd__o221a_1
X_5941_ _1023_ _1264_ VGND VGND VPWR VPWR 
+ _1802_
+ sky130_fd_sc_hd__or2_1
X_5942_ _1802_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__clkbuf_2
X_5943_ _1803_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__inv_2
X_5944_ \gpio_configure[5][12]\ _1803_ net359 _1804_ VGND VGND 
+ VPWR
+ VPWR _0347_ sky130_fd_sc_hd__a22o_1
X_5945_ \gpio_configure[5][11]\ _1803_ net361 _1804_ VGND VGND 
+ VPWR
+ VPWR _0346_ sky130_fd_sc_hd__a22o_1
X_5946_ \gpio_configure[5][10]\ _1803_ net363 _1804_ VGND VGND 
+ VPWR
+ VPWR _0345_ sky130_fd_sc_hd__a22o_1
X_5947_ \gpio_configure[5][9]\ _1803_ net366 _1804_ VGND VGND 
+ VPWR
+ VPWR _0344_ sky130_fd_sc_hd__a22o_1
X_5948_ \gpio_configure[5][8]\ _1803_ net367 _1804_ VGND VGND 
+ VPWR
+ VPWR _0343_ sky130_fd_sc_hd__a22o_1
X_5949_ _1022_ _1168_ VGND VGND VPWR VPWR 
+ _1805_
+ sky130_fd_sc_hd__or2_1
X_5950_ _1805_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__clkbuf_4
X_5951_ _1806_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__inv_2
X_5952_ \gpio_configure[4][7]\ _1806_ \cdata[7]\ _1807_ VGND VGND 
+ VPWR
+ VPWR _0342_ sky130_fd_sc_hd__a22o_1
X_5953_ \gpio_configure[4][6]\ _1806_ \cdata[6]\ _1807_ VGND VGND 
+ VPWR
+ VPWR _0341_ sky130_fd_sc_hd__a22o_1
X_5954_ \gpio_configure[4][5]\ _1806_ \cdata[5]\ _1807_ VGND VGND 
+ VPWR
+ VPWR _0340_ sky130_fd_sc_hd__a22o_1
X_5955_ \gpio_configure[4][4]\ _1806_ net360 _1807_ VGND VGND 
+ VPWR
+ VPWR _0339_ sky130_fd_sc_hd__a22o_1
X_5956_ \gpio_configure[4][3]\ _1806_ net362 _1807_ VGND VGND 
+ VPWR
+ VPWR _0338_ sky130_fd_sc_hd__a22o_1
X_5957_ \gpio_configure[4][2]\ _1806_ net364 _1807_ VGND VGND 
+ VPWR
+ VPWR _0337_ sky130_fd_sc_hd__a22o_1
X_5958_ \gpio_configure[4][1]\ _1806_ net366 _1807_ VGND VGND 
+ VPWR
+ VPWR _0336_ sky130_fd_sc_hd__a22o_1
X_5959_ \gpio_configure[4][0]\ _1806_ net368 _1807_ VGND VGND 
+ VPWR
+ VPWR _0335_ sky130_fd_sc_hd__a22o_1
X_5960_ _1023_ _1245_ VGND VGND VPWR VPWR 
+ _1808_
+ sky130_fd_sc_hd__or2_1
X_5961_ _1808_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__clkbuf_2
X_5962_ _1809_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__inv_2
X_5963_ \gpio_configure[4][12]\ _1809_ net359 _1810_ VGND VGND 
+ VPWR
+ VPWR _0334_ sky130_fd_sc_hd__a22o_1
X_5964_ \gpio_configure[4][11]\ _1809_ net361 _1810_ VGND VGND 
+ VPWR
+ VPWR _0333_ sky130_fd_sc_hd__a22o_1
X_5965_ \gpio_configure[4][10]\ _1809_ net363 _1810_ VGND VGND 
+ VPWR
+ VPWR _0332_ sky130_fd_sc_hd__a22o_1
X_5966_ \gpio_configure[4][9]\ _1809_ net365 _1810_ VGND VGND 
+ VPWR
+ VPWR _0331_ sky130_fd_sc_hd__a22o_1
X_5967_ \gpio_configure[4][8]\ _1809_ net367 _1810_ VGND VGND 
+ VPWR
+ VPWR _0330_ sky130_fd_sc_hd__a22o_1
X_5968_ _1022_ _1321_ VGND VGND VPWR VPWR 
+ _1811_
+ sky130_fd_sc_hd__or2_1
X_5969_ _1811_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__clkbuf_4
X_5970_ _1812_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__inv_2
X_5971_ \gpio_configure[3][7]\ _1812_ \cdata[7]\ _1813_ VGND VGND 
+ VPWR
+ VPWR _0329_ sky130_fd_sc_hd__a22o_1
X_5972_ \gpio_configure[3][6]\ _1812_ \cdata[6]\ _1813_ VGND VGND 
+ VPWR
+ VPWR _0328_ sky130_fd_sc_hd__a22o_1
X_5973_ \gpio_configure[3][5]\ _1812_ \cdata[5]\ _1813_ VGND VGND 
+ VPWR
+ VPWR _0327_ sky130_fd_sc_hd__a22o_1
X_5974_ \gpio_configure[3][4]\ _1812_ net360 _1813_ VGND VGND 
+ VPWR
+ VPWR _0326_ sky130_fd_sc_hd__a22o_1
X_5975_ \gpio_configure[3][3]\ _1812_ net362 _1813_ VGND VGND 
+ VPWR
+ VPWR _0325_ sky130_fd_sc_hd__a22o_1
X_5976_ \gpio_configure[3][2]\ _1812_ \cdata[2]\ _1813_ VGND VGND 
+ VPWR
+ VPWR _0324_ sky130_fd_sc_hd__a22o_1
X_5977_ \gpio_configure[3][1]\ _1812_ net366 _1813_ VGND VGND 
+ VPWR
+ VPWR _0323_ sky130_fd_sc_hd__a22o_1
X_5978_ \gpio_configure[3][0]\ _1812_ \cdata[0]\ _1813_ VGND VGND 
+ VPWR
+ VPWR _0322_ sky130_fd_sc_hd__a22o_1
X_5979_ _1449_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__clkbuf_1
X_5980_ _1814_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
X_5981_ \hkspi.count[0]\ _1465_ \hkspi.count[1]\ VGND VGND VPWR 
+ VPWR
+ _1815_ sky130_fd_sc_hd__and3_1
X_5982_ \hkspi.count[2]\ _1815_ _1419_ _1466_ VGND VGND 
+ VPWR
+ VPWR _0321_ sky130_fd_sc_hd__o22a_1
X_5983_ _1449_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__clkbuf_1
X_5984_ _1816_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_5985_ _1417_ _1466_ VGND VGND VPWR VPWR 
+ _1817_
+ sky130_fd_sc_hd__nor2_1
X_5986_ \hkspi.count[1]\ _1817_ _1815_ VGND VGND VPWR 
+ VPWR
+ _0320_ sky130_fd_sc_hd__o21ba_1
X_5987_ _1449_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__clkbuf_1
X_5988_ _1818_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
X_5989_ _1417_ _1466_ _1817_ VGND VGND VPWR 
+ VPWR
+ _0319_ sky130_fd_sc_hd__a21oi_1
X_5990_ _1449_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__clkbuf_1
X_5991_ _1819_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
X_5992_ \hkspi.fixed[0]\ _1442_ VGND VGND VPWR VPWR 
+ _1820_
+ sky130_fd_sc_hd__nand2_1
X_5993_ \hkspi.state[2]\ _1420_ _1820_ VGND VGND VPWR 
+ VPWR
+ _1821_ sky130_fd_sc_hd__and3_1
X_5994_ \hkspi.state[3]\ _1821_ _0087_ VGND VGND VPWR 
+ VPWR
+ _1822_ sky130_fd_sc_hd__o21ai_4
X_5995_ _1822_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__inv_2
X_5996_ \hkspi.addr[7]\ _1822_ _0054_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0318_ sky130_fd_sc_hd__a22o_1
X_5997_ _1449_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__clkbuf_1
X_5998_ _1824_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
X_5999_ \hkspi.addr[6]\ _1822_ _0053_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0317_ sky130_fd_sc_hd__a22o_1
X_6000_ _1449_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__clkbuf_1
X_6001_ _1825_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
X_6002_ \hkspi.addr[5]\ _1822_ _0052_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0316_ sky130_fd_sc_hd__a22o_1
X_6003_ _1449_ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__clkbuf_1
X_6004_ _1826_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
X_6005_ \hkspi.addr[4]\ _1822_ _0051_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0315_ sky130_fd_sc_hd__a22o_1
X_6006_ _1449_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__clkbuf_1
X_6007_ _1827_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
X_6008_ \hkspi.addr[3]\ _1822_ _0050_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0314_ sky130_fd_sc_hd__a22o_1
X_6009_ _1449_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__clkbuf_1
X_6010_ _1828_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
X_6011_ \hkspi.addr[2]\ _1822_ _0049_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0313_ sky130_fd_sc_hd__a22o_1
X_6012_ _1449_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__clkbuf_1
X_6013_ _1829_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
X_6014_ \hkspi.addr[1]\ _1822_ _0048_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0312_ sky130_fd_sc_hd__a22o_1
X_6015_ _1449_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__clkbuf_1
X_6016_ _1830_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
X_6017_ \hkspi.addr[0]\ _1822_ _0047_ _1823_ VGND VGND 
+ VPWR
+ VPWR _0311_ sky130_fd_sc_hd__a22o_1
X_6018_ net368 trap_output_dest _1048_ VGND VGND VPWR 
+ VPWR
+ _1831_ sky130_fd_sc_hd__mux2_1
X_6019_ _1831_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
X_6020_ _1449_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__clkbuf_1
X_6021_ _1832_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
X_6022_ _1415_ _0087_ _1417_ _1416_ VGND VGND 
+ VPWR
+ VPWR _1833_ sky130_fd_sc_hd__or4_1
X_6023_ _1833_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__inv_2
X_6024_ \hkspi.pre_pass_thru_user\ _1834_ \hkspi.pass_thru_user_delay\ _1833_ VGND VGND 
+ VPWR
+ VPWR _0309_ sky130_fd_sc_hd__a22o_1
X_6025_ serial_bb_data_1 _1034_ \cdata[5]\ _1035_ VGND VGND 
+ VPWR
+ VPWR _0308_ sky130_fd_sc_hd__a22o_1
X_6026_ serial_bb_resetn _1034_ net364 _1035_ VGND VGND 
+ VPWR
+ VPWR _0307_ sky130_fd_sc_hd__a22o_1
X_6027_ _1022_ _1293_ VGND VGND VPWR VPWR 
+ _1835_
+ sky130_fd_sc_hd__or2_1
X_6028_ _1835_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__clkbuf_4
X_6029_ _1836_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__inv_2
X_6030_ \gpio_configure[26][7]\ _1836_ \cdata[7]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0306_ sky130_fd_sc_hd__a22o_1
X_6031_ \gpio_configure[26][6]\ _1836_ \cdata[6]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0305_ sky130_fd_sc_hd__a22o_1
X_6032_ \gpio_configure[26][5]\ _1836_ \cdata[5]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0304_ sky130_fd_sc_hd__a22o_1
X_6033_ \gpio_configure[26][4]\ _1836_ \cdata[4]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0303_ sky130_fd_sc_hd__a22o_1
X_6034_ \gpio_configure[26][3]\ _1836_ \cdata[3]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0302_ sky130_fd_sc_hd__a22o_1
X_6035_ \gpio_configure[26][2]\ _1836_ \cdata[2]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0301_ sky130_fd_sc_hd__a22o_1
X_6036_ \gpio_configure[26][1]\ _1836_ \cdata[1]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0300_ sky130_fd_sc_hd__a22o_1
X_6037_ \gpio_configure[26][0]\ _1836_ \cdata[0]\ _1837_ VGND VGND 
+ VPWR
+ VPWR _0299_ sky130_fd_sc_hd__a22o_1
X_6038_ serial_bb_load _1034_ net362 _1035_ VGND VGND 
+ VPWR
+ VPWR _0298_ sky130_fd_sc_hd__a22o_1
X_6039__1 clknet_2_1_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR net379 sky130_fd_sc_hd__inv_4
X_6040_ _1449_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__clkbuf_1
X_6041_ _1838_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
X_6042_ _1126_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__clkbuf_1
X_6043_ _1839_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
X_6044_ _1126_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__clkbuf_1
X_6045_ _1840_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
X_6046_ _1126_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__clkbuf_1
X_6047_ _1841_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
X_6048_ _1126_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__clkbuf_1
X_6049_ _1842_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_1
X_6050_ _1126_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__clkbuf_1
X_6051_ _1843_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__clkbuf_1
X_6052_ _1022_ _1124_ _1161_ VGND VGND VPWR 
+ VPWR
+ _1844_ sky130_fd_sc_hd__or3_2
X_6053_ _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__clkbuf_2
X_6054_ _1845_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__inv_2
X_6055_ net303 _1845_ net362 _1846_ VGND VGND 
+ VPWR
+ VPWR _0297_ sky130_fd_sc_hd__a22o_1
X_6056_ net302 _1845_ net364 _1846_ VGND VGND 
+ VPWR
+ VPWR _0296_ sky130_fd_sc_hd__a22o_1
X_6057_ net301 _1845_ net366 _1846_ VGND VGND 
+ VPWR
+ VPWR _0295_ sky130_fd_sc_hd__a22o_1
X_6058_ net300 _1845_ net368 _1846_ VGND VGND 
+ VPWR
+ VPWR _0294_ sky130_fd_sc_hd__a22o_1
X_6059_ \gpio_configure[3][7]\ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__clkinv_2
X_6060_ net70 VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__inv_4
X_6061_ \gpio_configure[36][7]\ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__clkinv_2
X_6062_ \gpio_configure[1][7]\ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__inv_2
X_6063_ _1849_ _1251_ _1850_ _1249_ VGND VGND 
+ VPWR
+ VPWR _1851_ sky130_fd_sc_hd__o22a_1
X_6064_ _1847_ _1321_ _1848_ _1177_ _1851_ VGND 
+ VGND
+ VPWR VPWR _1852_ sky130_fd_sc_hd__o221a_1
X_6065_ \gpio_configure[8][7]\ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__clkinv_2
X_6066_ \gpio_configure[14][7]\ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__clkinv_2
X_6067_ \gpio_configure[37][7]\ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__inv_2
X_6068_ \gpio_configure[34][7]\ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__clkinv_2
X_6069_ _1855_ _1212_ _1856_ _1155_ VGND VGND 
+ VPWR
+ VPWR _1857_ sky130_fd_sc_hd__o22a_1
X_6070_ _1853_ _1196_ _1854_ _1206_ _1857_ VGND 
+ VGND
+ VPWR VPWR _1858_ sky130_fd_sc_hd__o221a_1
X_6071_ _1852_ _1858_ VGND VGND VPWR VPWR 
+ _1859_
+ sky130_fd_sc_hd__nand2_1
X_6072_ \gpio_configure[31][7]\ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__inv_2
X_6073_ \gpio_configure[29][7]\ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__inv_2
X_6074_ \gpio_configure[20][7]\ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__clkinv_4
X_6075_ net122 VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__clkinv_4
X_6076_ _1862_ _1392_ _1863_ _1339_ VGND VGND 
+ VPWR
+ VPWR _1864_ sky130_fd_sc_hd__o22a_1
X_6077_ _1860_ _1295_ _1861_ _1334_ _1864_ VGND 
+ VGND
+ VPWR VPWR _1865_ sky130_fd_sc_hd__o221a_1
X_6078_ \gpio_configure[22][7]\ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__clkinv_4
X_6079_ \gpio_configure[28][7]\ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__clkinv_2
X_6080_ \gpio_configure[33][7]\ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__clkinv_2
X_6081_ _1868_ _1224_ VGND VGND VPWR VPWR 
+ _1869_
+ sky130_fd_sc_hd__or2_1
X_6082_ _1866_ _1375_ _1867_ _1388_ _1869_ VGND 
+ VGND
+ VPWR VPWR _1870_ sky130_fd_sc_hd__o221a_2
X_6083_ \gpio_configure[27][7]\ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__clkinv_4
X_6084_ net297 VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__inv_2
X_6085_ net10 VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__inv_2
X_6086_ _1065_ _1167_ VGND VGND VPWR VPWR 
+ _1874_
+ sky130_fd_sc_hd__or2_4
X_6087_ net33 VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__inv_2
X_6088_ _1873_ _1874_ _1875_ _1348_ VGND VGND 
+ VPWR
+ VPWR _1876_ sky130_fd_sc_hd__o22a_1
X_6089_ _1871_ _1273_ _1872_ _1106_ _1876_ VGND 
+ VGND
+ VPWR VPWR _1877_ sky130_fd_sc_hd__o221a_2
X_6090_ \gpio_configure[19][7]\ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__inv_2
X_6091_ \gpio_configure[18][7]\ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__clkinv_2
X_6092_ net280 VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__inv_2
X_6093_ net19 VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__inv_2
X_6094_ _1880_ _1101_ _1881_ _1384_ VGND VGND 
+ VPWR
+ VPWR _1882_ sky130_fd_sc_hd__o22a_2
X_6095_ _1878_ _1406_ _1879_ _1355_ _1882_ VGND 
+ VGND
+ VPWR VPWR _1883_ sky130_fd_sc_hd__o221a_1
X_6096_ _1865_ _1870_ _1877_ _1883_ VGND VGND 
+ VPWR
+ VPWR _1884_ sky130_fd_sc_hd__and4_2
X_6097_ net117 VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__clkinv_2
X_6098_ \gpio_configure[17][7]\ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__inv_2
X_6099_ net99 VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__clkinv_2
X_6100_ net108 VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__inv_2
X_6101_ _1887_ _1370_ _1888_ _1319_ VGND VGND 
+ VPWR
+ VPWR _1889_ sky130_fd_sc_hd__o22a_1
X_6102_ _1885_ _1310_ _1886_ _1284_ _1889_ VGND 
+ VGND
+ VPWR VPWR _1890_ sky130_fd_sc_hd__o221a_2
X_6103_ \gpio_configure[32][7]\ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__clkinv_4
X_6104_ \gpio_configure[26][7]\ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__clkinv_4
X_6105_ \gpio_configure[0][7]\ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__inv_2
X_6106_ net28 VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__clkinv_2
X_6107_ _1893_ _1353_ _1894_ _1300_ VGND VGND 
+ VPWR
+ VPWR _1895_ sky130_fd_sc_hd__o22a_4
X_6108_ _1891_ _1312_ _1892_ _1293_ _1895_ VGND 
+ VGND
+ VPWR VPWR _1896_ sky130_fd_sc_hd__o221a_1
X_6109_ \gpio_configure[24][7]\ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__inv_2
X_6110_ \gpio_configure[23][7]\ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__inv_2
X_6111_ _1028_ _1070_ net323 VGND VGND VPWR 
+ VPWR
+ _1899_ sky130_fd_sc_hd__or3b_4
X_6112_ _1897_ _1325_ _1898_ _1404_ _1899_ VGND 
+ VGND
+ VPWR VPWR _1900_ sky130_fd_sc_hd__o221a_1
X_6113_ \gpio_configure[21][7]\ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__inv_2
X_6114_ \gpio_configure[30][7]\ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__clkinv_4
X_6115_ net289 VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__inv_2
X_6116_ \gpio_configure[25][7]\ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__inv_2
X_6117_ _1903_ _1096_ _1904_ _1054_ VGND VGND 
+ VPWR
+ VPWR _1905_ sky130_fd_sc_hd__o22a_2
X_6118_ _1901_ _1394_ _1902_ _1329_ _1905_ VGND 
+ VGND
+ VPWR VPWR _1906_ sky130_fd_sc_hd__o221a_1
X_6119_ _1890_ _1896_ _1900_ _1906_ VGND VGND 
+ VPWR
+ VPWR _1907_ sky130_fd_sc_hd__and4_1
X_6120_ \gpio_configure[5][7]\ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__clkinv_2
X_6121_ \gpio_configure[10][7]\ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__clkinv_2
X_6122_ \gpio_configure[12][7]\ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__inv_2
X_6123_ \gpio_configure[6][7]\ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__inv_2
X_6124_ _1910_ _1259_ _1911_ _1146_ VGND VGND 
+ VPWR
+ VPWR _1912_ sky130_fd_sc_hd__o22a_1
X_6125_ _1908_ _1181_ _1909_ _1214_ _1912_ VGND 
+ VGND
+ VPWR VPWR _1913_ sky130_fd_sc_hd__o221a_1
X_6126_ \gpio_configure[11][7]\ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__clkinv_2
X_6127_ \gpio_configure[4][7]\ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__inv_2
X_6128_ \gpio_configure[7][7]\ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__inv_2
X_6129_ \gpio_configure[2][7]\ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__clkinv_2
X_6130_ _1916_ _1149_ _1917_ _1253_ VGND VGND 
+ VPWR
+ VPWR _1918_ sky130_fd_sc_hd__o22a_1
X_6131_ _1914_ _1188_ _1915_ _1168_ _1918_ VGND 
+ VGND
+ VPWR VPWR _1919_ sky130_fd_sc_hd__o221a_1
X_6132_ net60 VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__inv_2
X_6133_ \gpio_configure[35][7]\ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__inv_2
X_6134_ _1218_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkinv_8
X_6135_ _1235_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkinv_8
X_6136_ net42 _0083_ net51 _0080_ VGND VGND 
+ VPWR
+ VPWR _1922_ sky130_fd_sc_hd__a22oi_1
X_6137_ _1920_ _1262_ _1921_ _1231_ _1922_ VGND 
+ VGND
+ VPWR VPWR _1923_ sky130_fd_sc_hd__o221a_2
X_6138_ \gpio_configure[15][7]\ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__clkinv_2
X_6139_ \gpio_configure[13][7]\ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__inv_2
X_6140_ \gpio_configure[9][7]\ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__inv_2
X_6141_ \gpio_configure[16][7]\ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__inv_2
X_6142_ _1926_ _1220_ _1927_ _1222_ VGND VGND 
+ VPWR
+ VPWR _1928_ sky130_fd_sc_hd__o22a_1
X_6143_ _1924_ _1239_ _1925_ _1200_ _1928_ VGND 
+ VGND
+ VPWR VPWR _1929_ sky130_fd_sc_hd__o221a_1
X_6144_ _1913_ _1919_ _1923_ _1929_ VGND VGND 
+ VPWR
+ VPWR _1930_ sky130_fd_sc_hd__and4_1
X_6145_ _1859_ _1884_ _1907_ _1930_ VGND VGND 
+ VPWR
+ VPWR \hkspi.idata[7]\ sky130_fd_sc_hd__nand4b_4
X_6146_ net196 VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__inv_2
X_6147_ _1931_ _1786_ VGND VGND VPWR VPWR 
+ _1932_
+ sky130_fd_sc_hd__or2_1
X_6148_ _1932_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__clkbuf_4
X_6149_ _1933_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__clkinv_2
X_6150_ \hkspi.idata[7]\ _1933_ net351 _1934_ VGND VGND 
+ VPWR
+ VPWR _0293_ sky130_fd_sc_hd__o22a_1
X_6151_ \gpio_configure[35][6]\ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__clkinv_2
X_6152_ \gpio_configure[18][6]\ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__inv_2
X_6153_ net32 VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__inv_2
X_6154_ \gpio_configure[17][6]\ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__clkinv_2
X_6155_ _1937_ _1348_ _1938_ _1284_ VGND VGND 
+ VPWR
+ VPWR _1939_ sky130_fd_sc_hd__o22a_1
X_6156_ _1935_ _1231_ _1936_ _1355_ _1939_ VGND 
+ VGND
+ VPWR VPWR _1940_ sky130_fd_sc_hd__o221a_1
X_6157_ \gpio_configure[1][6]\ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__inv_2
X_6158_ _1065_ _1114_ VGND VGND VPWR VPWR 
+ _1942_
+ sky130_fd_sc_hd__or2_4
X_6159_ \gpio_configure[21][6]\ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__inv_2
X_6160_ \gpio_configure[29][6]\ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__inv_2
X_6161_ _1943_ _1394_ _1944_ _1334_ VGND VGND 
+ VPWR
+ VPWR _1945_ sky130_fd_sc_hd__o22a_1
X_6162_ _1941_ _1249_ _1942_ _1945_ VGND VGND 
+ VPWR
+ VPWR _1946_ sky130_fd_sc_hd__o211a_1
X_6163_ \gpio_configure[36][6]\ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__inv_2
X_6164_ \gpio_configure[19][6]\ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__inv_2
X_6165_ _1177_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkinv_8
X_6166_ net69 _0085_ net50 _0080_ VGND VGND 
+ VPWR
+ VPWR _1949_ sky130_fd_sc_hd__a22oi_1
X_6167_ _1947_ _1251_ _1948_ _1406_ _1949_ VGND 
+ VGND
+ VPWR VPWR _1950_ sky130_fd_sc_hd__o221a_1
X_6168_ \gpio_configure[28][6]\ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__inv_2
X_6169_ \gpio_configure[23][6]\ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__inv_2
X_6170_ \gpio_configure[37][6]\ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__clkinv_2
X_6171_ \gpio_configure[24][6]\ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__inv_2
X_6172_ _1953_ _1212_ _1954_ _1325_ VGND VGND 
+ VPWR
+ VPWR _1955_ sky130_fd_sc_hd__o22a_1
X_6173_ _1951_ _1388_ _1952_ _1404_ _1955_ VGND 
+ VGND
+ VPWR VPWR _1956_ sky130_fd_sc_hd__o221a_1
X_6174_ _1940_ _1946_ _1950_ _1956_ VGND VGND 
+ VPWR
+ VPWR _1957_ sky130_fd_sc_hd__and4_1
X_6175_ \gpio_configure[9][6]\ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__clkinv_2
X_6176_ \gpio_configure[16][6]\ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__clkinv_2
X_6177_ _1958_ _1220_ _1959_ _1222_ VGND VGND 
+ VPWR
+ VPWR _1960_ sky130_fd_sc_hd__o22a_1
X_6178_ \gpio_configure[13][6]\ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__inv_2
X_6179_ \gpio_configure[14][6]\ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__clkinv_2
X_6180_ _1961_ _1200_ _1962_ _1206_ VGND VGND 
+ VPWR
+ VPWR _1963_ sky130_fd_sc_hd__o22a_1
X_6181_ \gpio_configure[15][6]\ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__inv_2
X_6182_ \gpio_configure[11][6]\ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__clkinv_2
X_6183_ \gpio_configure[12][6]\ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__clkinv_2
X_6184_ \gpio_configure[10][6]\ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__clkinv_2
X_6185_ _1966_ _1259_ _1967_ _1214_ VGND VGND 
+ VPWR
+ VPWR _1968_ sky130_fd_sc_hd__o22a_1
X_6186_ _1964_ _1239_ _1965_ _1188_ _1968_ VGND 
+ VGND
+ VPWR VPWR _1969_ sky130_fd_sc_hd__o221a_1
X_6187_ _1960_ _1963_ _1969_ VGND VGND VPWR 
+ VPWR
+ _1970_ sky130_fd_sc_hd__and3_1
X_6188_ \gpio_configure[26][6]\ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__clkinv_4
X_6189_ \gpio_configure[25][6]\ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__inv_2
X_6190_ \gpio_configure[32][6]\ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__clkinv_2
X_6191_ net41 _0083_ _1973_ _1312_ VGND VGND 
+ VPWR
+ VPWR _1974_ sky130_fd_sc_hd__o2bb2a_1
X_6192_ _1971_ _1293_ _1972_ _1054_ _1974_ VGND 
+ VGND
+ VPWR VPWR _1975_ sky130_fd_sc_hd__o221a_1
X_6193_ net59 VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__inv_2
X_6194_ \gpio_configure[8][6]\ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__clkinv_2
X_6195_ \gpio_configure[30][6]\ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__clkinv_2
X_6196_ \gpio_configure[22][6]\ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__inv_2
X_6197_ _1978_ _1329_ _1979_ _1375_ VGND VGND 
+ VPWR
+ VPWR _1980_ sky130_fd_sc_hd__o22a_1
X_6198_ _1976_ _1262_ _1977_ _1196_ _1980_ VGND 
+ VGND
+ VPWR VPWR _1981_ sky130_fd_sc_hd__o221a_1
X_6199_ \gpio_configure[27][6]\ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__inv_2
X_6200_ \gpio_configure[31][6]\ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__inv_2
X_6201_ \gpio_configure[33][6]\ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__clkinv_4
X_6202_ net296 VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__inv_2
X_6203_ _1984_ _1224_ _1985_ _1106_ VGND VGND 
+ VPWR
+ VPWR _1986_ sky130_fd_sc_hd__o22a_1
X_6204_ _1982_ _1273_ _1983_ _1295_ _1986_ VGND 
+ VGND
+ VPWR VPWR _1987_ sky130_fd_sc_hd__o221a_1
X_6205_ \gpio_configure[34][6]\ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__clkinv_4
X_6206_ net9 VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__inv_2
X_6207_ net27 VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__inv_2
X_6208_ net18 VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__inv_2
X_6209_ _1990_ _1300_ _1991_ _1384_ VGND VGND 
+ VPWR
+ VPWR _1992_ sky130_fd_sc_hd__o22a_1
X_6210_ _1988_ _1155_ _1989_ _1874_ _1992_ VGND 
+ VGND
+ VPWR VPWR _1993_ sky130_fd_sc_hd__o221a_2
X_6211_ _1975_ _1981_ _1987_ _1993_ VGND VGND 
+ VPWR
+ VPWR _1994_ sky130_fd_sc_hd__and4_1
X_6212_ \gpio_configure[7][6]\ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__clkinv_4
X_6213_ net308 VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__clkinv_2
X_6214_ net279 VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__clkinv_2
X_6215_ \gpio_configure[5][6]\ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__inv_2
X_6216_ _1997_ _1101_ _1998_ _1181_ VGND VGND 
+ VPWR
+ VPWR _1999_ sky130_fd_sc_hd__o22a_1
X_6217_ _1995_ _1149_ _1996_ _1032_ _1999_ VGND 
+ VGND
+ VPWR VPWR _2000_ sky130_fd_sc_hd__o221a_1
X_6218_ \gpio_configure[4][6]\ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__clkinv_4
X_6219_ net107 VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__clkinv_2
X_6220_ net288 VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__inv_2
X_6221_ net98 VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__clkinv_2
X_6222_ _2003_ _1096_ _2004_ _1370_ VGND VGND 
+ VPWR
+ VPWR _2005_ sky130_fd_sc_hd__o22a_1
X_6223_ _2001_ _1168_ _2002_ _1319_ _2005_ VGND 
+ VGND
+ VPWR VPWR _2006_ sky130_fd_sc_hd__o221a_1
X_6224_ \gpio_configure[6][6]\ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__clkinv_2
X_6225_ \gpio_configure[20][6]\ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__inv_2
X_6226_ net322 VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__clkinv_2
X_6227_ net116 VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__inv_2
X_6228_ _2009_ _1071_ _2010_ _1310_ VGND VGND 
+ VPWR
+ VPWR _2011_ sky130_fd_sc_hd__o22a_2
X_6229_ _2007_ _1146_ _2008_ _1392_ _2011_ VGND 
+ VGND
+ VPWR VPWR _2012_ sky130_fd_sc_hd__o221a_1
X_6230_ \gpio_configure[3][6]\ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__inv_2
X_6231_ \gpio_configure[0][6]\ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__inv_2
X_6232_ \gpio_configure[2][6]\ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__clkinv_2
X_6233_ net121 VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__clkinv_4
X_6234_ _2015_ _1253_ _2016_ _1339_ VGND VGND 
+ VPWR
+ VPWR _2017_ sky130_fd_sc_hd__o22a_1
X_6235_ _2013_ _1321_ _2014_ _1353_ _2017_ VGND 
+ VGND
+ VPWR VPWR _2018_ sky130_fd_sc_hd__o221a_1
X_6236_ _2000_ _2006_ _2012_ _2018_ VGND VGND 
+ VPWR
+ VPWR _2019_ sky130_fd_sc_hd__and4_2
X_6237_ _1957_ _1970_ _1994_ _2019_ VGND VGND 
+ VPWR
+ VPWR \hkspi.idata[6]\ sky130_fd_sc_hd__nand4_4
X_6238_ _1933_ \hkspi.idata[6]\ net350 _1934_ VGND VGND 
+ VPWR
+ VPWR _0292_ sky130_fd_sc_hd__o22a_1
X_6239_ \gpio_configure[20][5]\ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__inv_2
X_6240_ \gpio_configure[23][5]\ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__inv_2
X_6241_ \gpio_configure[25][5]\ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__inv_2
X_6242_ _2021_ _1404_ _2022_ _1054_ VGND VGND 
+ VPWR
+ VPWR _2023_ sky130_fd_sc_hd__o22a_1
X_6243_ net278 VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__inv_2
X_6244_ \gpio_configure[29][5]\ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__clkinv_4
X_6245_ net25 VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__clkinv_2
X_6246_ \gpio_configure[31][5]\ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__inv_2
X_6247_ _2026_ _1300_ _2027_ _1295_ VGND VGND 
+ VPWR
+ VPWR _2028_ sky130_fd_sc_hd__o22a_1
X_6248_ _2024_ _1101_ _2025_ _1334_ _2028_ VGND 
+ VGND
+ VPWR VPWR _2029_ sky130_fd_sc_hd__o221a_2
X_6249_ net114 VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__inv_2
X_6250_ \gpio_configure[0][5]\ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__inv_2
X_6251_ _1032_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__inv_4
X_6252_ net106 VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__clkinv_2
X_6253_ net307 _2032_ _2033_ _1319_ VGND VGND 
+ VPWR
+ VPWR _2034_ sky130_fd_sc_hd__o2bb2a_1
X_6254_ _2030_ _1310_ _2031_ _1353_ _2034_ VGND 
+ VGND
+ VPWR VPWR _2035_ sky130_fd_sc_hd__o221a_2
X_6255_ _2020_ _1392_ _2023_ _2029_ _2035_ VGND 
+ VGND
+ VPWR VPWR _2036_ sky130_fd_sc_hd__o2111a_1
X_6256_ \gpio_configure[30][5]\ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__inv_4
X_6257_ net31 VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__inv_2
X_6258_ net295 VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__inv_2
X_6259_ net8 VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__inv_2
X_6260_ _2039_ _1106_ _2040_ _1874_ VGND VGND 
+ VPWR
+ VPWR _2041_ sky130_fd_sc_hd__o22a_1
X_6261_ _2037_ _1329_ _2038_ _1348_ _2041_ VGND 
+ VGND
+ VPWR VPWR _2042_ sky130_fd_sc_hd__o221a_1
X_6262_ net17 VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__clkinv_2
X_6263_ \gpio_configure[27][5]\ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__clkinv_4
X_6264_ \gpio_configure[32][5]\ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__inv_6
X_6265_ net262 VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__inv_2
X_6266_ _2045_ _1312_ _2046_ _1110_ VGND VGND 
+ VPWR
+ VPWR _2047_ sky130_fd_sc_hd__o22a_1
X_6267_ _2043_ _1384_ _2044_ _1273_ _2047_ VGND 
+ VGND
+ VPWR VPWR _2048_ sky130_fd_sc_hd__o221a_1
X_6268_ net321 VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__clkinv_2
X_6269_ \gpio_configure[19][5]\ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__clkinv_4
X_6270_ net120 VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__clkinv_2
X_6271_ \gpio_configure[28][5]\ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__inv_6
X_6272_ _2051_ _1339_ _2052_ _1388_ VGND VGND 
+ VPWR
+ VPWR _2053_ sky130_fd_sc_hd__o22a_1
X_6273_ _2049_ _1071_ _2050_ _1406_ _2053_ VGND 
+ VGND
+ VPWR VPWR _2054_ sky130_fd_sc_hd__o221a_1
X_6274_ \gpio_configure[21][5]\ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__clkinv_4
X_6275_ \gpio_configure[24][5]\ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__inv_2
X_6276_ \gpio_configure[18][5]\ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__inv_2
X_6277_ \gpio_configure[17][5]\ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__inv_2
X_6278_ _2057_ _1355_ _2058_ _1284_ VGND VGND 
+ VPWR
+ VPWR _2059_ sky130_fd_sc_hd__o22a_1
X_6279_ _2055_ _1394_ _2056_ _1325_ _2059_ VGND 
+ VGND
+ VPWR VPWR _2060_ sky130_fd_sc_hd__o221a_2
X_6280_ _2042_ _2048_ _2054_ _2060_ VGND VGND 
+ VPWR
+ VPWR _2061_ sky130_fd_sc_hd__and4_2
X_6281_ net68 VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__inv_2
X_6282_ \gpio_configure[2][5]\ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__clkinv_2
X_6283_ \gpio_configure[15][5]\ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__clkinv_2
X_6284_ \gpio_configure[8][5]\ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__inv_2
X_6285_ _2064_ _1239_ _2065_ _1196_ VGND VGND 
+ VPWR
+ VPWR _2066_ sky130_fd_sc_hd__o22a_1
X_6286_ _2062_ _1177_ _2063_ _1253_ _2066_ VGND 
+ VGND
+ VPWR VPWR _2067_ sky130_fd_sc_hd__o221a_1
X_6287_ \gpio_configure[35][5]\ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__inv_2
X_6288_ \gpio_configure[10][5]\ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__inv_2
X_6289_ net287 VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__clkinv_2
X_6290_ \gpio_configure[22][5]\ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__inv_6
X_6291_ \gpio_configure[26][5]\ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__inv_6
X_6292_ net97 VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__clkinv_2
X_6293_ _2072_ _1293_ _2073_ _1370_ VGND VGND 
+ VPWR
+ VPWR _2074_ sky130_fd_sc_hd__o22a_1
X_6294_ _2070_ _1096_ _2071_ _1375_ _2074_ VGND 
+ VGND
+ VPWR VPWR _2075_ sky130_fd_sc_hd__o221a_4
X_6295_ _2068_ _1231_ _2069_ _1214_ _2075_ VGND 
+ VGND
+ VPWR VPWR _2076_ sky130_fd_sc_hd__o221a_1
X_6296_ \gpio_configure[37][5]\ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__inv_2
X_6297_ \gpio_configure[5][5]\ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__clkinv_2
X_6298_ \gpio_configure[9][5]\ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__inv_2
X_6299_ net49 _0080_ _2079_ _1220_ VGND VGND 
+ VPWR
+ VPWR _2080_ sky130_fd_sc_hd__o2bb2a_1
X_6300_ _2077_ _1212_ _2078_ _1181_ _2080_ VGND 
+ VGND
+ VPWR VPWR _2081_ sky130_fd_sc_hd__o221a_1
X_6301_ \gpio_configure[11][5]\ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__inv_2
X_6302_ \gpio_configure[7][5]\ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__clkinv_2
X_6303_ \gpio_configure[3][5]\ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__clkinv_2
X_6304_ \gpio_configure[6][5]\ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__inv_2
X_6305_ _2084_ _1321_ _2085_ _1146_ VGND VGND 
+ VPWR
+ VPWR _2086_ sky130_fd_sc_hd__o22a_1
X_6306_ _2082_ _1188_ _2083_ _1149_ _2086_ VGND 
+ VGND
+ VPWR VPWR _2087_ sky130_fd_sc_hd__o221a_1
X_6307_ _2067_ _2076_ _2081_ _2087_ VGND VGND 
+ VPWR
+ VPWR _2088_ sky130_fd_sc_hd__and4_1
X_6308_ \gpio_configure[12][5]\ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__clkinv_2
X_6309_ \gpio_configure[13][5]\ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__inv_2
X_6310_ \gpio_configure[33][5]\ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__clkinv_2
X_6311_ \gpio_configure[36][5]\ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__inv_2
X_6312_ _2091_ _1224_ _2092_ _1251_ VGND VGND 
+ VPWR
+ VPWR _2093_ sky130_fd_sc_hd__o22a_1
X_6313_ _2089_ _1259_ _2090_ _1200_ _2093_ VGND 
+ VGND
+ VPWR VPWR _2094_ sky130_fd_sc_hd__o221a_1
X_6314_ \gpio_configure[1][5]\ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__inv_2
X_6315_ \gpio_configure[4][5]\ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__clkinv_2
X_6316_ \gpio_configure[14][5]\ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__clkinv_2
X_6317_ net40 VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__inv_2
X_6318_ _2097_ _1206_ _2098_ _1218_ VGND VGND 
+ VPWR
+ VPWR _2099_ sky130_fd_sc_hd__o22a_1
X_6319_ _2095_ _1249_ _2096_ _1168_ _2099_ VGND 
+ VGND
+ VPWR VPWR _2100_ sky130_fd_sc_hd__o221a_1
X_6320_ \gpio_configure[16][5]\ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__clkinv_2
X_6321_ \gpio_configure[34][5]\ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__clkinv_2
X_6322_ _1262_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__inv_6
X_6323_ net66 _1159_ net57 _0081_ VGND VGND 
+ VPWR
+ VPWR _2103_ sky130_fd_sc_hd__a22oi_4
X_6324_ _2101_ _1222_ _2102_ _1155_ _2103_ VGND 
+ VGND
+ VPWR VPWR _2104_ sky130_fd_sc_hd__o221a_1
X_6325_ _2094_ _2100_ _2104_ VGND VGND VPWR 
+ VPWR
+ _2105_ sky130_fd_sc_hd__and3_2
X_6326_ _2036_ _2061_ _2088_ _2105_ VGND VGND 
+ VPWR
+ VPWR \hkspi.idata[5]\ sky130_fd_sc_hd__nand4_4
X_6327_ _1933_ \hkspi.idata[5]\ net348 _1934_ VGND VGND 
+ VPWR
+ VPWR _0291_ sky130_fd_sc_hd__o22a_1
X_6328_ \gpio_configure[19][4]\ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__clkinv_2
X_6329_ \gpio_configure[23][4]\ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__clkinv_4
X_6330_ \gpio_configure[24][12]\ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__clkinv_2
X_6331_ \gpio_configure[6][12]\ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__clkinv_2
X_6332_ _2108_ _1282_ _2109_ _1255_ VGND VGND 
+ VPWR
+ VPWR _2110_ sky130_fd_sc_hd__o22a_1
X_6333_ _2106_ _1406_ _2107_ _1404_ _2110_ VGND 
+ VGND
+ VPWR VPWR _2111_ sky130_fd_sc_hd__o221a_1
X_6334_ \gpio_configure[3][4]\ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__inv_2
X_6335_ \gpio_configure[34][12]\ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__inv_2
X_6336_ net96 VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__inv_2
X_6337_ \gpio_configure[6][4]\ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__clkinv_2
X_6338_ _2114_ _1370_ _2115_ _1146_ VGND VGND 
+ VPWR
+ VPWR _2116_ sky130_fd_sc_hd__o22a_1
X_6339_ _2112_ _1321_ _2113_ _1266_ _2116_ VGND 
+ VGND
+ VPWR VPWR _2117_ sky130_fd_sc_hd__o221a_1
X_6340_ \gpio_configure[28][12]\ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__clkinv_2
X_6341_ \gpio_configure[25][12]\ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__clkinv_2
X_6342_ net269 VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__clkinv_2
X_6343_ \gpio_configure[36][12]\ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__inv_2
X_6344_ _2120_ _1115_ _2121_ _1243_ VGND VGND 
+ VPWR
+ VPWR _2122_ sky130_fd_sc_hd__o22a_1
X_6345_ _2118_ _1361_ _2119_ _1288_ _2122_ VGND 
+ VGND
+ VPWR VPWR _2123_ sky130_fd_sc_hd__o221a_1
X_6346_ \gpio_configure[24][4]\ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__inv_2
X_6347_ \gpio_configure[23][12]\ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__clkinv_2
X_6348_ \gpio_configure[21][12]\ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__clkinv_2
X_6349_ \gpio_configure[28][4]\ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__clkinv_4
X_6350_ _2126_ _1377_ _2127_ _1388_ VGND VGND 
+ VPWR
+ VPWR _2128_ sky130_fd_sc_hd__o22a_1
X_6351_ _2124_ _1325_ _2125_ _1408_ _2128_ VGND 
+ VGND
+ VPWR VPWR _2129_ sky130_fd_sc_hd__o221a_1
X_6352_ _2111_ _2117_ _2123_ _2129_ VGND VGND 
+ VPWR
+ VPWR _2130_ sky130_fd_sc_hd__and4_1
X_6353_ \gpio_configure[9][4]\ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__clkinv_2
X_6354_ \gpio_configure[0][12]\ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__inv_2
X_6355_ _2132_ _1275_ _1322_ _1942_ VGND VGND 
+ VPWR
+ VPWR _2133_ sky130_fd_sc_hd__o211a_1
X_6356_ \gpio_configure[37][4]\ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__inv_2
X_6357_ \gpio_configure[20][4]\ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__inv_2
X_6358_ serial_bb_clock _2032_ _2135_ _1392_ VGND VGND 
+ VPWR
+ VPWR _2136_ sky130_fd_sc_hd__o2bb2a_2
X_6359_ net381 _1177_ _2134_ _1212_ _2136_ VGND 
+ VGND
+ VPWR VPWR _2137_ sky130_fd_sc_hd__o221a_2
X_6360_ \gpio_configure[16][4]\ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__clkinv_4
X_6361_ \gpio_configure[16][12]\ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__clkinv_2
X_6362_ \gpio_configure[13][12]\ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__inv_2
X_6363_ \gpio_configure[17][12]\ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__inv_2
X_6364_ _2140_ _1209_ _2141_ _1142_ VGND VGND 
+ VPWR
+ VPWR _2142_ sky130_fd_sc_hd__o22a_1
X_6365_ _2138_ _1222_ _2139_ _1198_ _2142_ VGND 
+ VGND
+ VPWR VPWR _2143_ sky130_fd_sc_hd__o221a_2
X_6366_ _2131_ _1220_ _2133_ _2137_ _2143_ VGND 
+ VGND
+ VPWR VPWR _2144_ sky130_fd_sc_hd__o2111a_2
X_6367_ \gpio_configure[10][4]\ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__clkinv_4
X_6368_ \gpio_configure[12][4]\ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__inv_2
X_6369_ \gpio_configure[10][12]\ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__inv_2
X_6370_ _2146_ _1259_ _2147_ _1165_ VGND VGND 
+ VPWR
+ VPWR _2148_ sky130_fd_sc_hd__o22a_1
X_6371_ \gpio_configure[13][4]\ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__inv_4
X_6372_ \gpio_configure[11][4]\ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__clkinv_2
X_6373_ \gpio_configure[11][12]\ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__clkinv_2
X_6374_ \gpio_configure[12][12]\ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__inv_2
X_6375_ _2151_ _1192_ _2152_ _1202_ VGND VGND 
+ VPWR
+ VPWR _2153_ sky130_fd_sc_hd__o22a_1
X_6376_ _2149_ _1200_ _2150_ _1188_ _2153_ VGND 
+ VGND
+ VPWR VPWR _2154_ sky130_fd_sc_hd__o221a_1
X_6377_ \gpio_configure[14][4]\ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__inv_2
X_6378_ \gpio_configure[15][12]\ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__clkinv_2
X_6379_ \gpio_configure[14][12]\ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__clkinv_2
X_6380_ \gpio_configure[15][4]\ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__inv_4
X_6381_ _2157_ _1186_ _2158_ _1239_ VGND VGND 
+ VPWR
+ VPWR _2159_ sky130_fd_sc_hd__o22a_1
X_6382_ _2155_ _1206_ _2156_ _1190_ _2159_ VGND 
+ VGND
+ VPWR VPWR _2160_ sky130_fd_sc_hd__o221a_2
X_6383_ _2145_ _1214_ _2148_ _2154_ _2160_ VGND 
+ VGND
+ VPWR VPWR _2161_ sky130_fd_sc_hd__o2111a_1
X_6384_ net286 VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__inv_2
X_6385_ net16 VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__inv_2
X_6386_ net7 VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__inv_2
X_6387_ \gpio_configure[30][12]\ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__clkinv_4
X_6388_ _2164_ _1874_ _2165_ _1344_ VGND VGND 
+ VPWR
+ VPWR _2166_ sky130_fd_sc_hd__o22a_1
X_6389_ _2162_ _1096_ _2163_ _1384_ _2166_ VGND 
+ VGND
+ VPWR VPWR _2167_ sky130_fd_sc_hd__o221a_2
X_6390_ \gpio_configure[30][4]\ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__clkinv_4
X_6391_ \gpio_configure[31][12]\ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__inv_2
X_6392_ \gpio_configure[33][4]\ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__inv_2
X_6393_ \gpio_configure[37][12]\ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__inv_2
X_6394_ _2170_ _1224_ _2171_ _1229_ VGND VGND 
+ VPWR
+ VPWR _2172_ sky130_fd_sc_hd__o22a_1
X_6395_ _2168_ _1329_ _2169_ _1337_ _2172_ VGND 
+ VGND
+ VPWR VPWR _2173_ sky130_fd_sc_hd__o221a_1
X_6396_ \gpio_configure[22][4]\ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__clkinv_4
X_6397_ \gpio_configure[29][12]\ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__inv_2
X_6398_ \gpio_configure[17][4]\ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__inv_2
X_6399_ \gpio_configure[22][12]\ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__inv_2
X_6400_ _2176_ _1284_ _2177_ _1402_ VGND VGND 
+ VPWR
+ VPWR _2178_ sky130_fd_sc_hd__o22a_1
X_6401_ _2174_ _1375_ _2175_ _1366_ _2178_ VGND 
+ VGND
+ VPWR VPWR _2179_ sky130_fd_sc_hd__o221a_1
X_6402_ \gpio_configure[27][4]\ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__inv_2
X_6403_ \gpio_configure[25][4]\ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__inv_2
X_6404_ \gpio_configure[19][12]\ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__clkinv_2
X_6405_ net277 VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__inv_2
X_6406_ _2182_ _1396_ _2183_ _1101_ VGND VGND 
+ VPWR
+ VPWR _2184_ sky130_fd_sc_hd__o22a_1
X_6407_ _2180_ _1273_ _2181_ _1054_ _2184_ VGND 
+ VGND
+ VPWR VPWR _2185_ sky130_fd_sc_hd__o221a_1
X_6408_ _2167_ _2173_ _2179_ _2185_ VGND VGND 
+ VPWR
+ VPWR _2186_ sky130_fd_sc_hd__and4_1
X_6409_ \gpio_configure[20][12]\ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__clkinv_2
X_6410_ \gpio_configure[36][4]\ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__clkinv_2
X_6411_ net24 VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__clkinv_2
X_6412_ \gpio_configure[27][12]\ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__inv_2
X_6413_ _2189_ _1300_ _2190_ _1315_ VGND VGND 
+ VPWR
+ VPWR _2191_ sky130_fd_sc_hd__o22a_2
X_6414_ _2187_ _1327_ _2188_ _1251_ _2191_ VGND 
+ VGND
+ VPWR VPWR _2192_ sky130_fd_sc_hd__o221a_1
X_6415_ \gpio_configure[21][4]\ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__clkinv_4
X_6416_ \gpio_configure[5][12]\ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__inv_2
X_6417_ \gpio_configure[32][12]\ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__inv_2
X_6418_ \gpio_configure[3][12]\ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__clkinv_4
X_6419_ _2195_ _1380_ _2196_ _1170_ VGND VGND 
+ VPWR
+ VPWR _2197_ sky130_fd_sc_hd__o22a_2
X_6420_ _2193_ _1394_ _2194_ _1264_ _2197_ VGND 
+ VGND
+ VPWR VPWR _2198_ sky130_fd_sc_hd__o221a_1
X_6421_ \gpio_configure[18][4]\ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__inv_2
X_6422_ \gpio_configure[31][4]\ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__clkinv_2
X_6423_ \gpio_configure[33][12]\ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__clkinv_2
X_6424_ \gpio_configure[18][12]\ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__inv_2
X_6425_ _2201_ _1368_ _2202_ _1398_ VGND VGND 
+ VPWR
+ VPWR _2203_ sky130_fd_sc_hd__o22a_1
X_6426_ _2199_ _1355_ _2200_ _1295_ _2203_ VGND 
+ VGND
+ VPWR VPWR _2204_ sky130_fd_sc_hd__o221a_1
X_6427_ \gpio_configure[29][4]\ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__clkinv_2
X_6428_ \gpio_configure[32][4]\ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__inv_2
X_6429_ \gpio_configure[26][12]\ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__clkinv_4
X_6430_ \gpio_configure[26][4]\ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__inv_4
X_6431_ _2207_ _1059_ _2208_ _1293_ VGND VGND 
+ VPWR
+ VPWR _2209_ sky130_fd_sc_hd__o22a_1
X_6432_ _2205_ _1334_ _2206_ _1312_ _2209_ VGND 
+ VGND
+ VPWR VPWR _2210_ sky130_fd_sc_hd__o221a_1
X_6433_ _2192_ _2198_ _2204_ _2210_ VGND VGND 
+ VPWR
+ VPWR _2211_ sky130_fd_sc_hd__and4_1
X_6434_ \gpio_configure[8][12]\ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__inv_2
X_6435_ \gpio_configure[0][4]\ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__inv_2
X_6436_ \gpio_configure[34][4]\ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__inv_2
X_6437_ _2213_ _1353_ _2214_ _1155_ VGND VGND 
+ VPWR
+ VPWR _2215_ sky130_fd_sc_hd__o22a_1
X_6438_ net105 VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__inv_2
X_6439_ \gpio_configure[1][4]\ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__clkinv_4
X_6440_ \gpio_configure[35][12]\ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__inv_2
X_6441_ \gpio_configure[7][12]\ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__clkinv_2
X_6442_ _2218_ _1151_ _2219_ _1179_ VGND VGND 
+ VPWR
+ VPWR _2220_ sky130_fd_sc_hd__o22a_1
X_6443_ _2216_ _1319_ _2217_ _1249_ _2220_ VGND 
+ VGND
+ VPWR VPWR _2221_ sky130_fd_sc_hd__o221a_1
X_6444_ net113 VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__inv_2
X_6445_ \gpio_configure[1][12]\ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__inv_2
X_6446_ net56 _0081_ net65 _1159_ VGND VGND 
+ VPWR
+ VPWR _2224_ sky130_fd_sc_hd__a22oi_4
X_6447_ _2222_ _1310_ _2223_ _1302_ _2224_ VGND 
+ VGND
+ VPWR VPWR _2225_ sky130_fd_sc_hd__o221a_1
X_6448_ _2212_ _1174_ _2215_ _2221_ _2225_ VGND 
+ VGND
+ VPWR VPWR _2226_ sky130_fd_sc_hd__o2111a_1
X_6449_ net294 VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__clkinv_2
X_6450_ net48 VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__clkinv_4
X_6451_ net119 VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__inv_2
X_6452_ net261 VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__inv_2
X_6453_ _2229_ _1339_ _2230_ _1110_ VGND VGND 
+ VPWR
+ VPWR _2231_ sky130_fd_sc_hd__o22a_2
X_6454_ _2227_ _1106_ _2228_ _1235_ _2231_ VGND 
+ VGND
+ VPWR VPWR _2232_ sky130_fd_sc_hd__o221a_1
X_6455_ net39 VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__clkinv_4
X_6456_ \gpio_configure[4][4]\ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__clkinv_2
X_6457_ \gpio_configure[8][4]\ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__inv_2
X_6458_ \gpio_configure[4][12]\ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__clkinv_4
X_6459_ _2235_ _1196_ _2236_ _1245_ VGND VGND 
+ VPWR
+ VPWR _2237_ sky130_fd_sc_hd__o22a_1
X_6460_ _2233_ _1218_ _2234_ _1168_ _2237_ VGND 
+ VGND
+ VPWR VPWR _2238_ sky130_fd_sc_hd__o221a_1
X_6461_ \gpio_configure[35][4]\ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__inv_2
X_6462_ \gpio_configure[5][4]\ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__clkinv_2
X_6463_ \gpio_configure[2][4]\ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__clkinv_2
X_6464_ \gpio_configure[2][12]\ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__inv_2
X_6465_ _2241_ _1253_ _2242_ _1157_ VGND VGND 
+ VPWR
+ VPWR _2243_ sky130_fd_sc_hd__o22a_1
X_6466_ _2239_ _1231_ _2240_ _1181_ _2243_ VGND 
+ VGND
+ VPWR VPWR _2244_ sky130_fd_sc_hd__o221a_1
X_6467_ \gpio_configure[9][12]\ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__inv_2
X_6468_ \gpio_configure[7][4]\ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__inv_2
X_6469_ net320 VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__inv_2
X_6470_ net30 VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__inv_2
X_6471_ _2247_ _1071_ _2248_ _1348_ VGND VGND 
+ VPWR
+ VPWR _2249_ sky130_fd_sc_hd__o22a_2
X_6472_ _2245_ _1241_ _2246_ _1149_ _2249_ VGND 
+ VGND
+ VPWR VPWR _2250_ sky130_fd_sc_hd__o221a_1
X_6473_ _2232_ _2238_ _2244_ _2250_ VGND VGND 
+ VPWR
+ VPWR _2251_ sky130_fd_sc_hd__and4_1
X_6474_ _2186_ _2211_ _2226_ _2251_ VGND VGND 
+ VPWR
+ VPWR _2252_ sky130_fd_sc_hd__and4_1
X_6475_ _2130_ _2144_ _2161_ _2252_ VGND VGND 
+ VPWR
+ VPWR \hkspi.idata[4]\ sky130_fd_sc_hd__nand4_2
X_6476_ _1933_ \hkspi.idata[4]\ net347 _1934_ VGND VGND 
+ VPWR
+ VPWR _0290_ sky130_fd_sc_hd__o22a_2
X_6477_ \gpio_configure[12][11]\ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__clkinv_2
X_6478_ \gpio_configure[13][3]\ VGND VGND VPWR VPWR _4419_ sky130_fd_sc_hd__inv_6
X_6479_ \gpio_configure[6][11]\ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__inv_2
X_6480_ \gpio_configure[36][11]\ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__inv_2
X_6481_ _2254_ _1255_ _2255_ _1243_ VGND VGND 
+ VPWR
+ VPWR _2256_ sky130_fd_sc_hd__o22a_1
X_6482_ _2253_ _1202_ _4419_ _1200_ _2256_ VGND 
+ VGND
+ VPWR VPWR _2257_ sky130_fd_sc_hd__o221a_1
X_6483_ \gpio_configure[15][3]\ VGND VGND VPWR VPWR _4421_ sky130_fd_sc_hd__inv_6
X_6484_ \gpio_configure[16][11]\ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__inv_2
X_6485_ \gpio_configure[36][3]\ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__inv_4
X_6486_ \gpio_configure[8][11]\ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__inv_2
X_6487_ _0093_ _1251_ _2259_ _1174_ VGND VGND 
+ VPWR
+ VPWR _2260_ sky130_fd_sc_hd__o22a_1
X_6488_ _4421_ _1239_ _2258_ _1198_ _2260_ VGND 
+ VGND
+ VPWR VPWR _2261_ sky130_fd_sc_hd__o221a_1
X_6489_ \gpio_configure[33][3]\ VGND VGND VPWR VPWR _4439_ sky130_fd_sc_hd__inv_4
X_6490_ \gpio_configure[3][3]\ VGND VGND VPWR VPWR _4409_ sky130_fd_sc_hd__inv_6
X_6491_ \gpio_configure[35][3]\ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__inv_2
X_6492_ \gpio_configure[10][3]\ VGND VGND VPWR VPWR _4416_ sky130_fd_sc_hd__inv_6
X_6493_ _0094_ _1231_ _4416_ _1214_ VGND VGND 
+ VPWR
+ VPWR _2262_ sky130_fd_sc_hd__o22a_1
X_6494_ _4439_ _1224_ _4409_ _1321_ _2262_ VGND 
+ VGND
+ VPWR VPWR _2263_ sky130_fd_sc_hd__o221a_2
X_6495_ \gpio_configure[15][11]\ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__inv_2
X_6496_ \gpio_configure[6][3]\ VGND VGND VPWR VPWR _4412_ sky130_fd_sc_hd__clkinv_4
X_6497_ \gpio_configure[13][11]\ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__clkinv_2
X_6498_ \gpio_configure[10][11]\ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__clkinv_2
X_6499_ _2265_ _1209_ _2266_ _1165_ VGND VGND 
+ VPWR
+ VPWR _2267_ sky130_fd_sc_hd__o22a_1
X_6500_ _2264_ _1190_ _4412_ _1146_ _2267_ VGND 
+ VGND
+ VPWR VPWR _2268_ sky130_fd_sc_hd__o221a_1
X_6501_ _2257_ _2261_ _2263_ _2268_ VGND VGND 
+ VPWR
+ VPWR _2269_ sky130_fd_sc_hd__and4_1
X_6502_ \gpio_configure[12][3]\ VGND VGND VPWR VPWR _4418_ sky130_fd_sc_hd__inv_6
X_6503_ \gpio_configure[34][11]\ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__inv_2
X_6504_ \gpio_configure[9][11]\ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__clkinv_4
X_6505_ net38 VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__inv_2
X_6506_ _2271_ _1241_ _2272_ _1218_ VGND VGND 
+ VPWR
+ VPWR _2273_ sky130_fd_sc_hd__o22a_1
X_6507_ _4418_ _1259_ _2270_ _1266_ _2273_ VGND 
+ VGND
+ VPWR VPWR _2274_ sky130_fd_sc_hd__o221a_1
X_6508_ \gpio_configure[17][11]\ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__inv_2
X_6509_ \gpio_configure[16][3]\ VGND VGND VPWR VPWR _4422_ sky130_fd_sc_hd__clkinv_8
X_6510_ \gpio_configure[14][11]\ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__inv_2
X_6511_ \gpio_configure[11][3]\ VGND VGND VPWR VPWR _4417_ sky130_fd_sc_hd__inv_6
X_6512_ _2276_ _1186_ _4417_ _1188_ VGND VGND 
+ VPWR
+ VPWR _2277_ sky130_fd_sc_hd__o22a_1
X_6513_ _2275_ _1142_ _4422_ _1222_ _2277_ VGND 
+ VGND
+ VPWR VPWR _2278_ sky130_fd_sc_hd__o221a_1
X_6514_ \gpio_configure[9][3]\ VGND VGND VPWR VPWR _4415_ sky130_fd_sc_hd__clkinv_4
X_6515_ \gpio_configure[14][3]\ VGND VGND VPWR VPWR _4420_ sky130_fd_sc_hd__inv_4
X_6516_ \gpio_configure[4][11]\ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__clkinv_4
X_6517_ \gpio_configure[1][3]\ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__inv_2
X_6518_ _2279_ _1245_ _2280_ _1249_ VGND VGND 
+ VPWR
+ VPWR _2281_ sky130_fd_sc_hd__o22a_1
X_6519_ _4415_ _1220_ _4420_ _1206_ _2281_ VGND 
+ VGND
+ VPWR VPWR _2282_ sky130_fd_sc_hd__o221a_1
X_6520_ \gpio_configure[8][3]\ VGND VGND VPWR VPWR _4414_ sky130_fd_sc_hd__clkinv_4
X_6521_ net46 VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__inv_4
X_6522_ \gpio_configure[37][11]\ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__clkinv_2
X_6523_ \gpio_configure[2][3]\ VGND VGND VPWR VPWR _4408_ sky130_fd_sc_hd__inv_4
X_6524_ _2284_ _1229_ _4408_ _1253_ VGND VGND 
+ VPWR
+ VPWR _2285_ sky130_fd_sc_hd__o22a_1
X_6525_ _4414_ _1196_ _2283_ _1235_ _2285_ VGND 
+ VGND
+ VPWR VPWR _2286_ sky130_fd_sc_hd__o221a_1
X_6526_ _2274_ _2278_ _2282_ _2286_ VGND VGND 
+ VPWR
+ VPWR _2287_ sky130_fd_sc_hd__and4_1
X_6527_ \gpio_configure[34][3]\ VGND VGND VPWR VPWR _4440_ sky130_fd_sc_hd__inv_6
X_6528_ \gpio_configure[7][11]\ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__inv_2
X_6529_ \gpio_configure[3][11]\ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__clkinv_4
X_6530_ _2288_ _1179_ _2289_ _1170_ VGND VGND 
+ VPWR
+ VPWR _2290_ sky130_fd_sc_hd__o22a_2
X_6531_ net55 VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__clkinv_4
X_6532_ \gpio_configure[7][3]\ VGND VGND VPWR VPWR _4413_ sky130_fd_sc_hd__clkinv_4
X_6533_ \gpio_configure[2][11]\ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__inv_2
X_6534_ net303 VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__inv_2
X_6535_ _2292_ _1157_ _2293_ _1161_ VGND VGND 
+ VPWR
+ VPWR _2294_ sky130_fd_sc_hd__o22a_1
X_6536_ _2291_ _1262_ _4413_ _1149_ _2294_ VGND 
+ VGND
+ VPWR VPWR _2295_ sky130_fd_sc_hd__o221a_1
X_6537_ \gpio_configure[4][3]\ VGND VGND VPWR VPWR _4410_ sky130_fd_sc_hd__clkinv_4
X_6538_ net64 VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__clkinv_4
X_6539_ \gpio_configure[5][11]\ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__inv_2
X_6540_ net67 _0085_ _2297_ _1264_ VGND VGND 
+ VPWR
+ VPWR _2298_ sky130_fd_sc_hd__o2bb2a_1
X_6541_ _4410_ _1168_ _2296_ _1158_ _2298_ VGND 
+ VGND
+ VPWR VPWR _2299_ sky130_fd_sc_hd__o221a_1
X_6542_ _4440_ _1155_ _2290_ _2295_ _2299_ VGND 
+ VGND
+ VPWR VPWR _2300_ sky130_fd_sc_hd__o2111a_1
X_6543_ \gpio_configure[31][11]\ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__clkinv_4
X_6544_ \gpio_configure[0][3]\ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkinv_2
X_6545_ net268 VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__inv_2
X_6546_ net276 VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__inv_2
X_6547_ _2302_ _1115_ _2303_ _1101_ VGND VGND 
+ VPWR
+ VPWR _2304_ sky130_fd_sc_hd__o22a_2
X_6548_ _2301_ _1337_ _0097_ _1353_ _2304_ VGND 
+ VGND
+ VPWR VPWR _2305_ sky130_fd_sc_hd__o221a_1
X_6549_ \gpio_configure[26][11]\ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__inv_2
X_6550_ \gpio_configure[28][11]\ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__inv_2
X_6551_ \gpio_configure[1][11]\ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__inv_2
X_6552_ net95 VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__inv_2
X_6553_ _2308_ _1302_ _2309_ _1370_ VGND VGND 
+ VPWR
+ VPWR _2310_ sky130_fd_sc_hd__o22a_1
X_6554_ _2306_ _1059_ _2307_ _1361_ _2310_ VGND 
+ VGND
+ VPWR VPWR _2311_ sky130_fd_sc_hd__o221a_1
X_6555_ \gpio_configure[18][11]\ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__clkinv_2
X_6556_ \gpio_configure[21][11]\ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__clkinv_2
X_6557_ \gpio_configure[33][11]\ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__inv_2
X_6558_ net103 VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__clkinv_2
X_6559_ _2314_ _1368_ _2315_ _1319_ VGND VGND 
+ VPWR
+ VPWR _2316_ sky130_fd_sc_hd__o22a_1
X_6560_ _2312_ _1398_ _2313_ _1377_ _2316_ VGND 
+ VGND
+ VPWR VPWR _2317_ sky130_fd_sc_hd__o221a_1
X_6561_ net112 VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__clkinv_2
X_6562_ \gpio_configure[30][3]\ VGND VGND VPWR VPWR _4436_ sky130_fd_sc_hd__inv_12
X_6563_ \gpio_configure[26][3]\ VGND VGND VPWR VPWR _4432_ sky130_fd_sc_hd__inv_8
X_6564_ net118 VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__inv_2
X_6565_ _4432_ _1293_ _2319_ _1339_ VGND VGND 
+ VPWR
+ VPWR _2320_ sky130_fd_sc_hd__o22a_1
X_6566_ _2318_ _1310_ _4436_ _1329_ _2320_ VGND 
+ VGND
+ VPWR VPWR _2321_ sky130_fd_sc_hd__o221a_1
X_6567_ _2305_ _2311_ _2317_ _2321_ VGND VGND 
+ VPWR
+ VPWR _2322_ sky130_fd_sc_hd__and4_1
X_6568_ \gpio_configure[29][3]\ VGND VGND VPWR VPWR _4435_ sky130_fd_sc_hd__clkinv_8
X_6569_ net293 VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__inv_2
X_6570_ net14 VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__clkinv_2
X_6571_ \gpio_configure[21][3]\ VGND VGND VPWR VPWR _4427_ sky130_fd_sc_hd__inv_6
X_6572_ _2324_ _1384_ _4427_ _1394_ VGND VGND 
+ VPWR
+ VPWR _2325_ sky130_fd_sc_hd__o22a_1
X_6573_ _4435_ _1334_ _2323_ _1106_ _2325_ VGND 
+ VGND
+ VPWR VPWR _2326_ sky130_fd_sc_hd__o221a_1
X_6574_ \gpio_configure[29][11]\ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__inv_2
X_6575_ \gpio_configure[18][3]\ VGND VGND VPWR VPWR _4424_ sky130_fd_sc_hd__clkinv_8
X_6576_ \gpio_configure[24][3]\ VGND VGND VPWR VPWR _4430_ sky130_fd_sc_hd__clkinv_8
X_6577_ \gpio_configure[32][11]\ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__inv_2
X_6578_ _4430_ _1325_ _2328_ _1380_ VGND VGND 
+ VPWR
+ VPWR _2329_ sky130_fd_sc_hd__o22a_1
X_6579_ _2327_ _1366_ _4424_ _1355_ _2329_ VGND 
+ VGND
+ VPWR VPWR _2330_ sky130_fd_sc_hd__o221a_1
X_6580_ \gpio_configure[5][3]\ VGND VGND VPWR VPWR _4411_ sky130_fd_sc_hd__clkinv_4
X_6581_ \gpio_configure[11][11]\ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__inv_2
X_6582_ \gpio_configure[37][3]\ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__inv_2
X_6583_ \gpio_configure[35][11]\ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__clkinv_4
X_6584_ _0092_ _1212_ _2332_ _1151_ VGND VGND 
+ VPWR
+ VPWR _2333_ sky130_fd_sc_hd__o22a_2
X_6585_ _4411_ _1181_ _2331_ _1192_ _2333_ VGND 
+ VGND
+ VPWR VPWR _2334_ sky130_fd_sc_hd__o221a_1
X_6586_ _2326_ _2330_ _2334_ VGND VGND VPWR 
+ VPWR
+ _2335_ sky130_fd_sc_hd__and3_1
X_6587_ \gpio_configure[19][11]\ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__inv_2
X_6588_ \gpio_configure[23][3]\ VGND VGND VPWR VPWR _4429_ sky130_fd_sc_hd__inv_6
X_6589_ \gpio_configure[22][11]\ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__inv_2
X_6590_ _4429_ _1404_ _2337_ _1402_ VGND VGND 
+ VPWR
+ VPWR _2338_ sky130_fd_sc_hd__o22a_2
X_6591_ net284 VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__inv_2
X_6592_ net6 VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__inv_2
X_6593_ net127 VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__clkinv_2
X_6594_ \gpio_configure[32][3]\ VGND VGND VPWR VPWR _4438_ sky130_fd_sc_hd__inv_6
X_6595_ _2341_ _1346_ _4438_ _1312_ VGND VGND 
+ VPWR
+ VPWR _2342_ sky130_fd_sc_hd__o22a_4
X_6596_ _2339_ _1096_ _2340_ _1874_ _2342_ VGND 
+ VGND
+ VPWR VPWR _2343_ sky130_fd_sc_hd__o221a_1
X_6597_ \gpio_configure[27][11]\ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__clkinv_2
X_6598_ \gpio_configure[27][3]\ VGND VGND VPWR VPWR _4433_ sky130_fd_sc_hd__inv_8
X_6599_ net260 VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__inv_2
X_6600_ serial_bb_load _2032_ _2345_ _1110_ VGND VGND 
+ VPWR
+ VPWR _2346_ sky130_fd_sc_hd__o2bb2a_1
X_6601_ _2344_ _1315_ _4433_ _1273_ _2346_ VGND 
+ VGND
+ VPWR VPWR _2347_ sky130_fd_sc_hd__o221a_1
X_6602_ _2336_ _1396_ _2338_ _2343_ _2347_ VGND 
+ VGND
+ VPWR VPWR _2348_ sky130_fd_sc_hd__o2111a_1
X_6603_ \gpio_configure[22][3]\ VGND VGND VPWR VPWR _4428_ sky130_fd_sc_hd__clkinv_8
X_6604_ \gpio_configure[23][11]\ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__clkinv_2
X_6605_ \gpio_configure[19][3]\ VGND VGND VPWR VPWR _4425_ sky130_fd_sc_hd__inv_8
X_6606_ \gpio_configure[24][11]\ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__clkinv_2
X_6607_ _4425_ _1406_ _2350_ _1282_ VGND VGND 
+ VPWR
+ VPWR _2351_ sky130_fd_sc_hd__o22a_1
X_6608_ _4428_ _1375_ _2349_ _1408_ _2351_ VGND 
+ VGND
+ VPWR VPWR _2352_ sky130_fd_sc_hd__o221a_1
X_6609_ \gpio_configure[25][11]\ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__clkinv_2
X_6610_ \gpio_configure[17][3]\ VGND VGND VPWR VPWR _4423_ sky130_fd_sc_hd__clkinv_8
X_6611_ \gpio_configure[20][3]\ VGND VGND VPWR VPWR _4426_ sky130_fd_sc_hd__inv_6
X_6612_ \gpio_configure[20][11]\ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__clkinv_2
X_6613_ _4426_ _1392_ _2354_ _1327_ VGND VGND 
+ VPWR
+ VPWR _2355_ sky130_fd_sc_hd__o22a_1
X_6614_ _2353_ _1288_ _4423_ _1284_ _2355_ VGND 
+ VGND
+ VPWR VPWR _2356_ sky130_fd_sc_hd__o221a_1
X_6615_ \gpio_configure[30][11]\ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__clkinv_4
X_6616_ \gpio_configure[31][3]\ VGND VGND VPWR VPWR _4437_ sky130_fd_sc_hd__clkinv_8
X_6617_ \gpio_configure[0][11]\ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__inv_2
X_6618_ net29 VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__inv_2
X_6619_ _2358_ _1275_ _2359_ _1348_ VGND VGND 
+ VPWR
+ VPWR _2360_ sky130_fd_sc_hd__o22a_1
X_6620_ _2357_ _1344_ _4437_ _1295_ _2360_ VGND 
+ VGND
+ VPWR VPWR _2361_ sky130_fd_sc_hd__o221a_1
X_6621_ net319 VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__clkinv_2
X_6622_ \gpio_configure[28][3]\ VGND VGND VPWR VPWR _4434_ sky130_fd_sc_hd__inv_8
X_6623_ \gpio_configure[25][3]\ VGND VGND VPWR VPWR _4431_ sky130_fd_sc_hd__inv_6
X_6624_ net23 VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__clkinv_2
X_6625_ _4431_ _1054_ _2363_ _1300_ VGND VGND 
+ VPWR
+ VPWR _2364_ sky130_fd_sc_hd__o22a_1
X_6626_ _2362_ _1071_ _4434_ _1388_ _2364_ VGND 
+ VGND
+ VPWR VPWR _2365_ sky130_fd_sc_hd__o221a_1
X_6627_ _2352_ _2356_ _2361_ _2365_ VGND VGND 
+ VPWR
+ VPWR _2366_ sky130_fd_sc_hd__and4_1
X_6628_ _2322_ _2335_ _2348_ _2366_ VGND VGND 
+ VPWR
+ VPWR _2367_ sky130_fd_sc_hd__and4_2
X_6629_ _2269_ _2287_ _2300_ _2367_ VGND VGND 
+ VPWR
+ VPWR \hkspi.idata[3]\ sky130_fd_sc_hd__nand4_4
X_6630_ _1933_ \hkspi.idata[3]\ net346 _1934_ VGND VGND 
+ VPWR
+ VPWR _0289_ sky130_fd_sc_hd__o22a_1
X_6631_ \gpio_configure[15][2]\ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__inv_2
X_6632_ \gpio_configure[16][10]\ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__clkinv_2
X_6633_ \gpio_configure[14][2]\ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__clkinv_2
X_6634_ \gpio_configure[14][10]\ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__clkinv_2
X_6635_ _2370_ _1206_ _2371_ _1186_ VGND VGND 
+ VPWR
+ VPWR _2372_ sky130_fd_sc_hd__o22a_1
X_6636_ _2368_ _1239_ _2369_ _1198_ _2372_ VGND 
+ VGND
+ VPWR VPWR _2373_ sky130_fd_sc_hd__o221a_1
X_6637_ \gpio_configure[10][2]\ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__inv_2
X_6638_ \gpio_configure[12][10]\ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__clkinv_2
X_6639_ \gpio_configure[11][2]\ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__clkinv_2
X_6640_ \gpio_configure[11][10]\ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__clkinv_2
X_6641_ _2376_ _1188_ _2377_ _1192_ VGND VGND 
+ VPWR
+ VPWR _2378_ sky130_fd_sc_hd__o22a_1
X_6642_ _2374_ _1214_ _2375_ _1202_ _2378_ VGND 
+ VGND
+ VPWR VPWR _2379_ sky130_fd_sc_hd__o221a_1
X_6643_ \gpio_configure[12][2]\ VGND VGND VPWR VPWR _2380_ sky130_fd_sc_hd__clkinv_2
X_6644_ \gpio_configure[9][2]\ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__inv_2
X_6645_ \gpio_configure[13][10]\ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__clkinv_2
X_6646_ \gpio_configure[10][10]\ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__inv_2
X_6647_ _2382_ _1209_ _2383_ _1165_ VGND VGND 
+ VPWR
+ VPWR _2384_ sky130_fd_sc_hd__o22a_1
X_6648_ _2380_ _1259_ _2381_ _1220_ _2384_ VGND 
+ VGND
+ VPWR VPWR _2385_ sky130_fd_sc_hd__o221a_1
X_6649_ _2373_ _2379_ _2385_ VGND VGND VPWR 
+ VPWR
+ _2386_ sky130_fd_sc_hd__and3_1
X_6650_ \gpio_configure[26][2]\ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__inv_4
X_6651_ net273 VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__inv_2
X_6652_ \gpio_configure[26][10]\ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__clkinv_4
X_6653_ net63 VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__inv_2
X_6654_ _2389_ _1059_ _2390_ _1158_ VGND VGND 
+ VPWR
+ VPWR _2391_ sky130_fd_sc_hd__o22a_1
X_6655_ _2387_ _1293_ _2388_ _1110_ _2391_ VGND 
+ VGND
+ VPWR VPWR _2392_ sky130_fd_sc_hd__o221a_1
X_6656_ net318 VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__inv_2
X_6657_ \gpio_configure[32][10]\ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__inv_2
X_6658_ clk1_output_dest VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__clkinv_4
X_6659_ _1058_ _1065_ _2395_ _1047_ _1942_ VGND 
+ VGND
+ VPWR VPWR _2396_ sky130_fd_sc_hd__o221a_1
X_6660_ _2393_ _1071_ _2394_ _1380_ _2396_ VGND 
+ VGND
+ VPWR VPWR _2397_ sky130_fd_sc_hd__o221a_1
X_6661_ \gpio_configure[16][2]\ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__clkinv_2
X_6662_ \gpio_configure[17][10]\ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__clkinv_2
X_6663_ \gpio_configure[15][10]\ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__inv_2
X_6664_ \gpio_configure[13][2]\ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__clkinv_4
X_6665_ _2400_ _1190_ _2401_ _1200_ VGND VGND 
+ VPWR
+ VPWR _2402_ sky130_fd_sc_hd__o22a_1
X_6666_ _2398_ _1222_ _2399_ _1142_ _2402_ VGND 
+ VGND
+ VPWR VPWR _2403_ sky130_fd_sc_hd__o221a_1
X_6667_ \gpio_configure[2][2]\ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__inv_2
X_6668_ \gpio_configure[34][10]\ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__inv_2
X_6669_ net111 VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__inv_2
X_6670_ net292 VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__clkinv_2
X_6671_ _2406_ _1310_ _2407_ _1106_ VGND VGND 
+ VPWR
+ VPWR _2408_ sky130_fd_sc_hd__o22a_1
X_6672_ _2404_ _1253_ _2405_ _1266_ _2408_ VGND 
+ VGND
+ VPWR VPWR _2409_ sky130_fd_sc_hd__o221a_1
X_6673_ \gpio_configure[3][2]\ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__clkinv_2
X_6674_ \gpio_configure[8][10]\ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__inv_2
X_6675_ net267 VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__inv_2
X_6676_ net129 VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__inv_4
X_6677_ _2412_ _1115_ _2413_ _1346_ VGND VGND 
+ VPWR
+ VPWR _2414_ sky130_fd_sc_hd__o22a_2
X_6678_ _2410_ _1321_ _2411_ _1174_ _2414_ VGND 
+ VGND
+ VPWR VPWR _2415_ sky130_fd_sc_hd__o221a_1
X_6679_ net115 VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__inv_4
X_6680_ net54 VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__clkinv_4
X_6681_ \gpio_configure[5][2]\ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__inv_2
X_6682_ \gpio_configure[9][10]\ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__clkinv_4
X_6683_ _2418_ _1181_ _2419_ _1241_ VGND VGND 
+ VPWR
+ VPWR _2420_ sky130_fd_sc_hd__o22a_1
X_6684_ _2416_ _1339_ _2417_ _1262_ _2420_ VGND 
+ VGND
+ VPWR VPWR _2421_ sky130_fd_sc_hd__o221a_1
X_6685_ \gpio_configure[3][10]\ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__clkinv_4
X_6686_ \gpio_configure[34][2]\ VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__inv_2
X_6687_ \gpio_configure[8][2]\ VGND VGND VPWR VPWR _2424_ sky130_fd_sc_hd__clkinv_2
X_6688_ net45 _0080_ _2424_ _1196_ VGND VGND 
+ VPWR
+ VPWR _2425_ sky130_fd_sc_hd__o2bb2a_1
X_6689_ _2422_ _1170_ _2423_ _1155_ _2425_ VGND 
+ VGND
+ VPWR VPWR _2426_ sky130_fd_sc_hd__o221a_1
X_6690_ _2409_ _2415_ _2421_ _2426_ VGND VGND 
+ VPWR
+ VPWR _2427_ sky130_fd_sc_hd__and4_1
X_6691_ _2392_ _2397_ _2403_ _2427_ VGND VGND 
+ VPWR
+ VPWR _2428_ sky130_fd_sc_hd__and4_1
X_6692_ \gpio_configure[25][2]\ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__inv_2
X_6693_ \gpio_configure[35][2]\ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__clkinv_2
X_6694_ \gpio_configure[24][2]\ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__inv_2
X_6695_ \gpio_configure[20][10]\ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__clkinv_2
X_6696_ _2431_ _1325_ _2432_ _1327_ VGND VGND 
+ VPWR
+ VPWR _2433_ sky130_fd_sc_hd__o22a_1
X_6697_ _2429_ _1054_ _2430_ _1231_ _2433_ VGND 
+ VGND
+ VPWR VPWR _2434_ sky130_fd_sc_hd__o221a_1
X_6698_ serial_bb_resetn VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__clkinv_2
X_6699_ net275 VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__inv_2
X_6700_ \gpio_configure[19][10]\ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__inv_2
X_6701_ \gpio_configure[36][10]\ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__inv_2
X_6702_ _2437_ _1396_ _2438_ _1243_ VGND VGND 
+ VPWR
+ VPWR _2439_ sky130_fd_sc_hd__o22a_2
X_6703_ _2435_ _1032_ _2436_ _1101_ _2439_ VGND 
+ VGND
+ VPWR VPWR _2440_ sky130_fd_sc_hd__o221a_4
X_6704_ \gpio_configure[30][2]\ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__inv_2
X_6705_ \gpio_configure[30][10]\ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__clkinv_4
X_6706_ net26 VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__clkinv_4
X_6707_ \gpio_configure[37][10]\ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__inv_2
X_6708_ _2443_ _1348_ _2444_ _1229_ VGND VGND 
+ VPWR
+ VPWR _2445_ sky130_fd_sc_hd__o22a_1
X_6709_ _2441_ _1329_ _2442_ _1344_ _2445_ VGND 
+ VGND
+ VPWR VPWR _2446_ sky130_fd_sc_hd__o221a_1
X_6710_ \gpio_configure[20][2]\ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__inv_2
X_6711_ \gpio_configure[28][10]\ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__clkinv_4
X_6712_ \gpio_configure[31][10]\ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__inv_2
X_6713_ \gpio_configure[21][2]\ VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__inv_2
X_6714_ _2449_ _1337_ _2450_ _1394_ VGND VGND 
+ VPWR
+ VPWR _2451_ sky130_fd_sc_hd__o22a_1
X_6715_ _2447_ _1392_ _2448_ _1361_ _2451_ VGND 
+ VGND
+ VPWR VPWR _2452_ sky130_fd_sc_hd__o221a_1
X_6716_ _2434_ _2440_ _2446_ _2452_ VGND VGND 
+ VPWR
+ VPWR _2453_ sky130_fd_sc_hd__and4_1
X_6717_ \gpio_configure[29][2]\ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__clkinv_2
X_6718_ \gpio_configure[18][10]\ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__inv_2
X_6719_ \gpio_configure[33][10]\ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__clkinv_2
X_6720_ \gpio_configure[32][2]\ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__inv_2
X_6721_ _2456_ _1368_ _2457_ _1312_ VGND VGND 
+ VPWR
+ VPWR _2458_ sky130_fd_sc_hd__o22a_1
X_6722_ _2454_ _1334_ _2455_ _1398_ _2458_ VGND 
+ VGND
+ VPWR VPWR _2459_ sky130_fd_sc_hd__o221a_1
X_6723_ \gpio_configure[21][10]\ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__inv_2
X_6724_ \gpio_configure[18][2]\ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__clkinv_2
X_6725_ \gpio_configure[27][10]\ VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__clkinv_2
X_6726_ net22 VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__clkinv_2
X_6727_ _2462_ _1315_ _2463_ _1300_ VGND VGND 
+ VPWR
+ VPWR _2464_ sky130_fd_sc_hd__o22a_2
X_6728_ _2460_ _1377_ _2461_ _1355_ _2464_ VGND 
+ VGND
+ VPWR VPWR _2465_ sky130_fd_sc_hd__o221a_1
X_6729_ \gpio_configure[22][10]\ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__clkinv_2
X_6730_ \gpio_configure[29][10]\ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__clkinv_2
X_6731_ \gpio_configure[4][10]\ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__clkinv_2
X_6732_ \gpio_configure[2][10]\ VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__inv_2
X_6733_ _2468_ _1245_ _2469_ _1157_ VGND VGND 
+ VPWR
+ VPWR _2470_ sky130_fd_sc_hd__o22a_1
X_6734_ _2466_ _1402_ _2467_ _1366_ _2470_ VGND 
+ VGND
+ VPWR VPWR _2471_ sky130_fd_sc_hd__o221a_1
X_6735_ \gpio_configure[28][2]\ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__clkinv_2
X_6736_ \gpio_configure[22][2]\ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__clkinv_4
X_6737_ \gpio_configure[17][2]\ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__inv_2
X_6738_ \gpio_configure[36][2]\ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__inv_2
X_6739_ _2474_ _1284_ _2475_ _1251_ VGND VGND 
+ VPWR
+ VPWR _2476_ sky130_fd_sc_hd__o22a_1
X_6740_ _2472_ _1388_ _2473_ _1375_ _2476_ VGND 
+ VGND
+ VPWR VPWR _2477_ sky130_fd_sc_hd__o221a_1
X_6741_ _2459_ _2465_ _2471_ _2477_ VGND VGND 
+ VPWR
+ VPWR _2478_ sky130_fd_sc_hd__and4_1
X_6742_ \gpio_configure[0][2]\ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__inv_2
X_6743_ \gpio_configure[6][10]\ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__clkinv_2
X_6744_ net102 VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__inv_2
X_6745_ \gpio_configure[1][10]\ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__clkinv_4
X_6746_ _2481_ _1319_ _2482_ _1302_ VGND VGND 
+ VPWR
+ VPWR _2483_ sky130_fd_sc_hd__o22a_1
X_6747_ _2479_ _1353_ _2480_ _1255_ _2483_ VGND 
+ VGND
+ VPWR VPWR _2484_ sky130_fd_sc_hd__o221a_2
X_6748_ \gpio_configure[37][2]\ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__inv_2
X_6749_ net302 VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__clkinv_4
X_6750_ \gpio_configure[7][10]\ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__inv_2
X_6751_ net37 _0083_ _2487_ _1179_ VGND VGND 
+ VPWR
+ VPWR _2488_ sky130_fd_sc_hd__o2bb2a_1
X_6752_ _2485_ _1212_ _2486_ _1161_ _2488_ VGND 
+ VGND
+ VPWR VPWR _2489_ sky130_fd_sc_hd__o221a_1
X_6753_ \gpio_configure[33][2]\ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__inv_2
X_6754_ \gpio_configure[6][2]\ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__clkinv_2
X_6755_ \gpio_configure[7][2]\ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__inv_2
X_6756_ \gpio_configure[35][10]\ VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__clkinv_2
X_6757_ _2492_ _1149_ _2493_ _1151_ VGND VGND 
+ VPWR
+ VPWR _2494_ sky130_fd_sc_hd__o22a_1
X_6758_ _2490_ _1224_ _2491_ _1146_ _2494_ VGND 
+ VGND
+ VPWR VPWR _2495_ sky130_fd_sc_hd__o221a_1
X_6759_ _2484_ _2489_ _2495_ VGND VGND VPWR 
+ VPWR
+ _2496_ sky130_fd_sc_hd__and3_1
X_6760_ \gpio_configure[23][2]\ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__clkinv_4
X_6761_ \gpio_configure[27][2]\ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__inv_2
X_6762_ \gpio_configure[25][10]\ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__clkinv_2
X_6763_ \gpio_configure[31][2]\ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__inv_2
X_6764_ _2499_ _1288_ _2500_ _1295_ VGND VGND 
+ VPWR
+ VPWR _2501_ sky130_fd_sc_hd__o22a_1
X_6765_ _2497_ _1404_ _2498_ _1273_ _2501_ VGND 
+ VGND
+ VPWR VPWR _2502_ sky130_fd_sc_hd__o221a_1
X_6766_ net13 VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__inv_2
X_6767_ \gpio_configure[19][2]\ VGND VGND VPWR VPWR _2504_ sky130_fd_sc_hd__clkinv_4
X_6768_ net283 VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__inv_2
X_6769_ net5 VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__inv_2
X_6770_ _2505_ _1096_ _2506_ _1874_ VGND VGND 
+ VPWR
+ VPWR _2507_ sky130_fd_sc_hd__o22a_1
X_6771_ _2503_ _1384_ _2504_ _1406_ _2507_ VGND 
+ VGND
+ VPWR VPWR _2508_ sky130_fd_sc_hd__o221a_1
X_6772_ \gpio_configure[5][10]\ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__inv_2
X_6773_ \gpio_configure[1][2]\ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__inv_2
X_6774_ \gpio_configure[0][10]\ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__inv_2
X_6775_ \gpio_configure[4][2]\ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__clkinv_4
X_6776_ _2511_ _1275_ _2512_ _1168_ VGND VGND 
+ VPWR
+ VPWR _2513_ sky130_fd_sc_hd__o22a_1
X_6777_ _2509_ _1264_ _2510_ _1249_ _2513_ VGND 
+ VGND
+ VPWR VPWR _2514_ sky130_fd_sc_hd__o221a_1
X_6778_ net94 VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__inv_2
X_6779_ \gpio_configure[24][10]\ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__inv_2
X_6780_ \gpio_configure[23][10]\ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__clkinv_2
X_6781_ _2516_ _1282_ _2517_ _1408_ VGND VGND 
+ VPWR
+ VPWR _2518_ sky130_fd_sc_hd__o22a_1
X_6782_ _2515_ _1370_ _1422_ _1177_ _2518_ VGND 
+ VGND
+ VPWR VPWR _2519_ sky130_fd_sc_hd__o221a_1
X_6783_ _2502_ _2508_ _2514_ _2519_ VGND VGND 
+ VPWR
+ VPWR _2520_ sky130_fd_sc_hd__and4_2
X_6784_ _2453_ _2478_ _2496_ _2520_ VGND VGND 
+ VPWR
+ VPWR _2521_ sky130_fd_sc_hd__and4_1
X_6785_ _2386_ _2428_ _2521_ VGND VGND VPWR 
+ VPWR
+ \hkspi.idata[2]\ sky130_fd_sc_hd__nand3_4
X_6786_ _1933_ \hkspi.idata[2]\ net345 _1934_ VGND VGND 
+ VPWR
+ VPWR _0288_ sky130_fd_sc_hd__o22a_1
X_6787_ \gpio_configure[30][1]\ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__clkinv_4
X_6788_ \gpio_configure[24][1]\ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__inv_2
X_6789_ net272 VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__inv_2
X_6790_ net317 VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__inv_2
X_6791_ _2524_ _1110_ _2525_ _1071_ VGND VGND 
+ VPWR
+ VPWR _2526_ sky130_fd_sc_hd__o22a_4
X_6792_ _2522_ _1329_ _2523_ _1325_ _2526_ VGND 
+ VGND
+ VPWR VPWR _2527_ sky130_fd_sc_hd__o221a_1
X_6793_ \gpio_configure[17][1]\ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__clkinv_4
X_6794_ net12 VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__inv_2
X_6795_ net324 VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__inv_2
X_6796_ net282 VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__inv_2
X_6797_ _2530_ _1076_ _2531_ _1096_ VGND VGND 
+ VPWR
+ VPWR _2532_ sky130_fd_sc_hd__o22a_2
X_6798_ _2528_ _1284_ _2529_ _1384_ _2532_ VGND 
+ VGND
+ VPWR VPWR _2533_ sky130_fd_sc_hd__o221a_1
X_6799_ \gpio_configure[6][1]\ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__inv_2
X_6800_ \gpio_configure[5][9]\ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__inv_2
X_6801_ \gpio_configure[18][9]\ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__inv_2
X_6802_ \gpio_configure[37][9]\ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__clkinv_2
X_6803_ _2536_ _1398_ _2537_ _1229_ _1942_ VGND 
+ VGND
+ VPWR VPWR _2538_ sky130_fd_sc_hd__o221a_1
X_6804_ _2534_ _1146_ _2535_ _1264_ _2538_ VGND 
+ VGND
+ VPWR VPWR _2539_ sky130_fd_sc_hd__o221a_1
X_6805_ \gpio_configure[27][9]\ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__clkinv_2
X_6806_ net101 VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__clkinv_2
X_6807_ clk2_output_dest VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__inv_4
X_6808_ net124 VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__clkinv_2
X_6809_ _2542_ _1047_ _2543_ _1370_ VGND VGND 
+ VPWR
+ VPWR _2544_ sky130_fd_sc_hd__o22a_1
X_6810_ _2540_ _1315_ _2541_ _1319_ _2544_ VGND 
+ VGND
+ VPWR VPWR _2545_ sky130_fd_sc_hd__o221a_1
X_6811_ net266 VGND VGND VPWR VPWR _2546_ sky130_fd_sc_hd__inv_2
X_6812_ \gpio_configure[26][9]\ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__clkinv_4
X_6813_ net15 VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__inv_2
X_6814_ net264 VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__inv_2
X_6815_ _2548_ _1348_ _2549_ _1120_ VGND VGND 
+ VPWR
+ VPWR _2550_ sky130_fd_sc_hd__o22a_1
X_6816_ _2546_ _1115_ _2547_ _1059_ _2550_ VGND 
+ VGND
+ VPWR VPWR _2551_ sky130_fd_sc_hd__o221a_1
X_6817_ net110 VGND VGND VPWR VPWR _2552_ sky130_fd_sc_hd__clkinv_2
X_6818_ \gpio_configure[31][1]\ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__clkinv_4
X_6819_ \gpio_configure[32][1]\ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__inv_4
X_6820_ net104 VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__inv_2
X_6821_ _2554_ _1312_ _2555_ _1339_ VGND VGND 
+ VPWR
+ VPWR _2556_ sky130_fd_sc_hd__o22a_1
X_6822_ _2552_ _1310_ _2553_ _1295_ _2556_ VGND 
+ VGND
+ VPWR VPWR _2557_ sky130_fd_sc_hd__o221a_1
X_6823_ \gpio_configure[26][1]\ VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__clkinv_4
X_6824_ \gpio_configure[30][9]\ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__inv_2
X_6825_ \gpio_configure[29][1]\ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__clkinv_2
X_6826_ \gpio_configure[32][9]\ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__inv_2
X_6827_ _2560_ _1334_ _2561_ _1380_ VGND VGND 
+ VPWR
+ VPWR _2562_ sky130_fd_sc_hd__o22a_1
X_6828_ _2558_ _1293_ _2559_ _1344_ _2562_ VGND 
+ VGND
+ VPWR VPWR _2563_ sky130_fd_sc_hd__o221a_2
X_6829_ _2545_ _2551_ _2557_ _2563_ VGND VGND 
+ VPWR
+ VPWR _2564_ sky130_fd_sc_hd__and4_1
X_6830_ _2527_ _2533_ _2539_ _2564_ VGND VGND 
+ VPWR
+ VPWR _2565_ sky130_fd_sc_hd__and4_1
X_6831_ net21 VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__clkinv_2
X_6832_ \gpio_configure[28][1]\ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__inv_6
X_6833_ \gpio_configure[1][9]\ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__clkinv_2
X_6834_ net285 VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__inv_2
X_6835_ _2568_ _1302_ _2569_ _1106_ VGND VGND 
+ VPWR
+ VPWR _2570_ sky130_fd_sc_hd__o22a_1
X_6836_ _2566_ _1300_ _2567_ _1388_ _2570_ VGND 
+ VGND
+ VPWR VPWR _2571_ sky130_fd_sc_hd__o221a_1
X_6837_ \gpio_configure[0][9]\ VGND VGND VPWR VPWR _2572_ sky130_fd_sc_hd__inv_2
X_6838_ \gpio_configure[0][1]\ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__inv_2
X_6839_ net291 VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__inv_2
X_6840_ \gpio_configure[33][9]\ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__inv_2
X_6841_ _2574_ _1092_ _2575_ _1368_ VGND VGND 
+ VPWR
+ VPWR _2576_ sky130_fd_sc_hd__o22a_1
X_6842_ _2572_ _1275_ _2573_ _1353_ _2576_ VGND 
+ VGND
+ VPWR VPWR _2577_ sky130_fd_sc_hd__o221a_1
X_6843_ \gpio_configure[23][9]\ VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__clkinv_2
X_6844_ \gpio_configure[25][1]\ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__inv_2
X_6845_ \gpio_configure[28][9]\ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__inv_2
X_6846_ _2579_ _1054_ _2580_ _1361_ VGND VGND 
+ VPWR
+ VPWR _2581_ sky130_fd_sc_hd__o22a_1
X_6847_ net128 VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__inv_4
X_6848_ \gpio_configure[29][9]\ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__clkinv_2
X_6849_ net35 VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__inv_2
X_6850_ serial_bb_enable _2032_ _2584_ _1874_ VGND VGND 
+ VPWR
+ VPWR _2585_ sky130_fd_sc_hd__o2bb2a_2
X_6851_ _2582_ _1346_ _2583_ _1366_ _2585_ VGND 
+ VGND
+ VPWR VPWR _2586_ sky130_fd_sc_hd__o221a_1
X_6852_ _2578_ _1408_ _2581_ _2586_ VGND VGND 
+ VPWR
+ VPWR _2587_ sky130_fd_sc_hd__o211a_1
X_6853_ \gpio_configure[21][1]\ VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__inv_2
X_6854_ \gpio_configure[23][1]\ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__inv_2
X_6855_ \gpio_configure[20][1]\ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__clkinv_2
X_6856_ \gpio_configure[31][9]\ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__clkinv_2
X_6857_ _2590_ _1392_ _2591_ _1337_ VGND VGND 
+ VPWR
+ VPWR _2592_ sky130_fd_sc_hd__o22a_1
X_6858_ _2588_ _1394_ _2589_ _1404_ _2592_ VGND 
+ VGND
+ VPWR VPWR _2593_ sky130_fd_sc_hd__o221a_2
X_6859_ \gpio_configure[18][1]\ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__inv_2
X_6860_ \gpio_configure[27][1]\ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__inv_2
X_6861_ net299 VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__inv_2
X_6862_ irq_2_inputsrc VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__clkinv_2
X_6863_ _2596_ _1101_ _2597_ _1304_ VGND VGND 
+ VPWR
+ VPWR _2598_ sky130_fd_sc_hd__o22a_2
X_6864_ _2594_ _1355_ _2595_ _1273_ _2598_ VGND 
+ VGND
+ VPWR VPWR _2599_ sky130_fd_sc_hd__o221a_1
X_6865_ \gpio_configure[22][1]\ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__inv_4
X_6866_ \gpio_configure[22][9]\ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__clkinv_2
X_6867_ \gpio_configure[20][9]\ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__clkinv_2
X_6868_ \gpio_configure[25][9]\ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__inv_2
X_6869_ _2602_ _1327_ _2603_ _1288_ VGND VGND 
+ VPWR
+ VPWR _2604_ sky130_fd_sc_hd__o22a_1
X_6870_ _2600_ _1375_ _2601_ _1402_ _2604_ VGND 
+ VGND
+ VPWR VPWR _2605_ sky130_fd_sc_hd__o221a_1
X_6871_ \gpio_configure[19][1]\ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__clkinv_4
X_6872_ \gpio_configure[19][9]\ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__clkinv_2
X_6873_ \gpio_configure[21][9]\ VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__clkinv_2
X_6874_ \gpio_configure[24][9]\ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__inv_2
X_6875_ _2608_ _1377_ _2609_ _1282_ VGND VGND 
+ VPWR
+ VPWR _2610_ sky130_fd_sc_hd__o22a_1
X_6876_ _2606_ _1406_ _2607_ _1396_ _2610_ VGND 
+ VGND
+ VPWR VPWR _2611_ sky130_fd_sc_hd__o221a_1
X_6877_ _2593_ _2599_ _2605_ _2611_ VGND VGND 
+ VPWR
+ VPWR _2612_ sky130_fd_sc_hd__and4_1
X_6878_ _2571_ _2577_ _2587_ _2612_ VGND VGND 
+ VPWR
+ VPWR _2613_ sky130_fd_sc_hd__and4_1
X_6879_ \gpio_configure[10][1]\ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__inv_2
X_6880_ \gpio_configure[15][1]\ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__inv_2
X_6881_ net47 _0085_ net53 _0081_ VGND VGND 
+ VPWR
+ VPWR _2616_ sky130_fd_sc_hd__a22oi_1
X_6882_ _2614_ _1214_ _2615_ _1239_ _2616_ VGND 
+ VGND
+ VPWR VPWR _2617_ sky130_fd_sc_hd__o221a_1
X_6883_ \gpio_configure[9][9]\ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__inv_2
X_6884_ \gpio_configure[36][1]\ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__clkinv_2
X_6885_ \gpio_configure[36][9]\ VGND VGND VPWR VPWR _2620_ sky130_fd_sc_hd__inv_2
X_6886_ net301 VGND VGND VPWR VPWR _2621_ sky130_fd_sc_hd__inv_2
X_6887_ _2620_ _1243_ _2621_ _1161_ VGND VGND 
+ VPWR
+ VPWR _2622_ sky130_fd_sc_hd__o22a_1
X_6888_ _2618_ _1241_ _2619_ _1251_ _2622_ VGND 
+ VGND
+ VPWR VPWR _2623_ sky130_fd_sc_hd__o221a_1
X_6889_ \gpio_configure[7][1]\ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__clkinv_2
X_6890_ \gpio_configure[11][1]\ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__clkinv_2
X_6891_ \gpio_configure[13][1]\ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__clkinv_4
X_6892_ \gpio_configure[34][9]\ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__clkinv_2
X_6893_ _2626_ _1200_ _2627_ _1266_ VGND VGND 
+ VPWR
+ VPWR _2628_ sky130_fd_sc_hd__o22a_1
X_6894_ _2624_ _1149_ _2625_ _1188_ _2628_ VGND 
+ VGND
+ VPWR VPWR _2629_ sky130_fd_sc_hd__o221a_1
X_6895_ \gpio_configure[16][1]\ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__clkinv_2
X_6896_ \gpio_configure[7][9]\ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__clkinv_2
X_6897_ \gpio_configure[10][9]\ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__clkinv_2
X_6898_ \gpio_configure[17][9]\ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__inv_2
X_6899_ _2632_ _1165_ _2633_ _1142_ VGND VGND 
+ VPWR
+ VPWR _2634_ sky130_fd_sc_hd__o22a_1
X_6900_ _2630_ _1222_ _2631_ _1179_ _2634_ VGND 
+ VGND
+ VPWR VPWR _2635_ sky130_fd_sc_hd__o221a_1
X_6901_ _2617_ _2623_ _2629_ _2635_ VGND VGND 
+ VPWR
+ VPWR _2636_ sky130_fd_sc_hd__and4_1
X_6902_ \gpio_configure[3][9]\ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__inv_4
X_6903_ net44 VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__inv_2
X_6904_ \gpio_configure[35][9]\ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__clkinv_4
X_6905_ \gpio_configure[33][1]\ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__clkinv_2
X_6906_ _2639_ _1151_ _2640_ _1224_ VGND VGND 
+ VPWR
+ VPWR _2641_ sky130_fd_sc_hd__o22a_1
X_6907_ _2637_ _1170_ _2638_ _1235_ _2641_ VGND 
+ VGND
+ VPWR VPWR _2642_ sky130_fd_sc_hd__o221a_1
X_6908_ \gpio_configure[1][1]\ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__inv_2
X_6909_ \gpio_configure[8][9]\ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__clkinv_4
X_6910_ \gpio_configure[2][1]\ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__inv_2
X_6911_ net62 _1159_ _2645_ _1253_ VGND VGND 
+ VPWR
+ VPWR _2646_ sky130_fd_sc_hd__o2bb2a_1
X_6912_ _2643_ _1249_ _2644_ _1174_ _2646_ VGND 
+ VGND
+ VPWR VPWR _2647_ sky130_fd_sc_hd__o221a_1
X_6913_ \gpio_configure[3][1]\ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__clkinv_2
X_6914_ \gpio_configure[37][1]\ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__clkinv_2
X_6915_ \gpio_configure[34][1]\ VGND VGND VPWR VPWR _2650_ sky130_fd_sc_hd__clkinv_2
X_6916_ \gpio_configure[35][1]\ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__inv_2
X_6917_ _2650_ _1155_ _2651_ _1231_ VGND VGND 
+ VPWR
+ VPWR _2652_ sky130_fd_sc_hd__o22a_1
X_6918_ _2648_ _1321_ _2649_ _1212_ _2652_ VGND 
+ VGND
+ VPWR VPWR _2653_ sky130_fd_sc_hd__o221a_1
X_6919_ \gpio_configure[4][1]\ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__clkinv_2
X_6920_ \gpio_configure[8][1]\ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__clkinv_2
X_6921_ \gpio_configure[5][1]\ VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__inv_2
X_6922_ \gpio_configure[6][9]\ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__clkinv_2
X_6923_ _2656_ _1181_ _2657_ _1255_ VGND VGND 
+ VPWR
+ VPWR _2658_ sky130_fd_sc_hd__o22a_1
X_6924_ _2654_ _1168_ _2655_ _1196_ _2658_ VGND 
+ VGND
+ VPWR VPWR _2659_ sky130_fd_sc_hd__o221a_1
X_6925_ _2642_ _2647_ _2653_ _2659_ VGND VGND 
+ VPWR
+ VPWR _2660_ sky130_fd_sc_hd__and4_1
X_6926_ \gpio_configure[14][1]\ VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__inv_2
X_6927_ \gpio_configure[13][9]\ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__inv_2
X_6928_ \gpio_configure[14][9]\ VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__clkinv_2
X_6929_ \gpio_configure[4][9]\ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__inv_2
X_6930_ _2663_ _1186_ _2664_ _1245_ VGND VGND 
+ VPWR
+ VPWR _2665_ sky130_fd_sc_hd__o22a_1
X_6931_ _2661_ _1206_ _2662_ _1209_ _2665_ VGND 
+ VGND
+ VPWR VPWR _2666_ sky130_fd_sc_hd__o221a_1
X_6932_ \gpio_configure[11][9]\ VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__inv_2
X_6933_ \gpio_configure[9][1]\ VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__inv_2
X_6934_ \gpio_configure[15][9]\ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__clkinv_2
X_6935_ \gpio_configure[12][9]\ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__inv_2
X_6936_ _2669_ _1190_ _2670_ _1202_ VGND VGND 
+ VPWR
+ VPWR _2671_ sky130_fd_sc_hd__o22a_1
X_6937_ _2667_ _1192_ _2668_ _1220_ _2671_ VGND 
+ VGND
+ VPWR VPWR _2672_ sky130_fd_sc_hd__o221a_1
X_6938_ \gpio_configure[16][9]\ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__clkinv_2
X_6939_ \gpio_configure[12][1]\ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__clkinv_2
X_6940_ \gpio_configure[2][9]\ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__clkinv_2
X_6941_ net72 VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__inv_2
X_6942_ _2675_ _1157_ _2676_ _1218_ VGND VGND 
+ VPWR
+ VPWR _2677_ sky130_fd_sc_hd__o22a_1
X_6943_ _2673_ _1198_ _2674_ _1259_ _2677_ VGND 
+ VGND
+ VPWR VPWR _2678_ sky130_fd_sc_hd__o221a_1
X_6944_ _2666_ _2672_ _2678_ VGND VGND VPWR 
+ VPWR
+ _2679_ sky130_fd_sc_hd__and3_1
X_6945_ _2636_ _2660_ _2679_ VGND VGND VPWR 
+ VPWR
+ _2680_ sky130_fd_sc_hd__and3_2
X_6946_ _2565_ _2613_ _2680_ VGND VGND VPWR 
+ VPWR
+ \hkspi.idata[1]\ sky130_fd_sc_hd__nand3_4
X_6947_ _1933_ \hkspi.idata[1]\ net344 _1934_ VGND VGND 
+ VPWR
+ VPWR _0287_ sky130_fd_sc_hd__o22a_1
X_6948_ _1413_ _1933_ net343 _1934_ VGND VGND 
+ VPWR
+ VPWR _0286_ sky130_fd_sc_hd__o22a_1
X_6949_ \wbbd_state[4]\ VGND VGND VPWR VPWR _2681_ sky130_fd_sc_hd__inv_2
X_6950_ _1931_ _2681_ VGND VGND VPWR VPWR 
+ _2682_
+ sky130_fd_sc_hd__or2_1
X_6951_ _2682_ VGND VGND VPWR VPWR _2683_ sky130_fd_sc_hd__clkbuf_4
X_6952_ _2683_ VGND VGND VPWR VPWR _2684_ sky130_fd_sc_hd__clkinv_2
X_6953_ \hkspi.idata[7]\ _2683_ net342 _2684_ VGND VGND 
+ VPWR
+ VPWR _0285_ sky130_fd_sc_hd__o22a_1
X_6954_ \hkspi.idata[6]\ _2683_ net341 _2684_ VGND VGND 
+ VPWR
+ VPWR _0284_ sky130_fd_sc_hd__o22a_1
X_6955_ \hkspi.idata[5]\ _2683_ net340 _2684_ VGND VGND 
+ VPWR
+ VPWR _0283_ sky130_fd_sc_hd__o22a_1
X_6956_ \hkspi.idata[4]\ _2683_ net339 _2684_ VGND VGND 
+ VPWR
+ VPWR _0282_ sky130_fd_sc_hd__o22a_2
X_6957_ \hkspi.idata[3]\ _2683_ net337 _2684_ VGND VGND 
+ VPWR
+ VPWR _0281_ sky130_fd_sc_hd__o22a_1
X_6958_ \hkspi.idata[2]\ _2683_ net336 _2684_ VGND VGND 
+ VPWR
+ VPWR _0280_ sky130_fd_sc_hd__o22a_1
X_6959_ \hkspi.idata[1]\ _2683_ net335 _2684_ VGND VGND 
+ VPWR
+ VPWR _0279_ sky130_fd_sc_hd__o22a_1
X_6960_ _1413_ _2683_ net334 _2684_ VGND VGND 
+ VPWR
+ VPWR _0278_ sky130_fd_sc_hd__o22a_1
X_6961_ \wbbd_state[3]\ VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__inv_2
X_6962_ _1931_ _2685_ VGND VGND VPWR VPWR 
+ _2686_
+ sky130_fd_sc_hd__or2_2
X_6963_ _2686_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__clkbuf_4
X_6964_ _2687_ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__inv_2
X_6965_ \hkspi.idata[7]\ _2687_ net356 _2688_ VGND VGND 
+ VPWR
+ VPWR _0277_ sky130_fd_sc_hd__o22a_1
X_6966_ \hkspi.idata[6]\ _2687_ net355 _2688_ VGND VGND 
+ VPWR
+ VPWR _0276_ sky130_fd_sc_hd__o22a_1
X_6967_ \hkspi.idata[5]\ _2687_ net354 _2688_ VGND VGND 
+ VPWR
+ VPWR _0275_ sky130_fd_sc_hd__o22a_1
X_6968_ \hkspi.idata[4]\ _2687_ net353 _2688_ VGND VGND 
+ VPWR
+ VPWR _0274_ sky130_fd_sc_hd__o22a_2
X_6969_ \hkspi.idata[3]\ _2687_ net352 _2688_ VGND VGND 
+ VPWR
+ VPWR _0273_ sky130_fd_sc_hd__o22a_1
X_6970_ \hkspi.idata[2]\ _2687_ net349 _2688_ VGND VGND 
+ VPWR
+ VPWR _0272_ sky130_fd_sc_hd__o22a_1
X_6971_ \hkspi.idata[1]\ _2687_ net338 _2688_ VGND VGND 
+ VPWR
+ VPWR _0271_ sky130_fd_sc_hd__o22a_1
X_6972_ _1413_ _2687_ net327 _2688_ VGND VGND 
+ VPWR
+ VPWR _0270_ sky130_fd_sc_hd__o22a_1
X_6973_ \wbbd_state[2]\ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__inv_2
X_6974_ _2689_ _1931_ VGND VGND VPWR VPWR 
+ _2690_
+ sky130_fd_sc_hd__or2_1
X_6975_ _2690_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__clkbuf_4
X_6976_ _2691_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__clkinv_2
X_6977_ \hkspi.idata[7]\ _2691_ net333 _2692_ VGND VGND 
+ VPWR
+ VPWR _0269_ sky130_fd_sc_hd__o22a_1
X_6978_ \hkspi.idata[6]\ _2691_ net332 _2692_ VGND VGND 
+ VPWR
+ VPWR _0268_ sky130_fd_sc_hd__o22a_1
X_6979_ \hkspi.idata[5]\ _2691_ net331 _2692_ VGND VGND 
+ VPWR
+ VPWR _0267_ sky130_fd_sc_hd__o22a_1
X_6980_ \hkspi.idata[4]\ _2691_ net330 _2692_ VGND VGND 
+ VPWR
+ VPWR _0266_ sky130_fd_sc_hd__o22a_2
X_6981_ \hkspi.idata[3]\ _2691_ net329 _2692_ VGND VGND 
+ VPWR
+ VPWR _0265_ sky130_fd_sc_hd__o22a_1
X_6982_ \hkspi.idata[2]\ _2691_ net328 _2692_ VGND VGND 
+ VPWR
+ VPWR _0264_ sky130_fd_sc_hd__o22a_1
X_6983_ \hkspi.idata[1]\ _2691_ net358 _2692_ VGND VGND 
+ VPWR
+ VPWR _0263_ sky130_fd_sc_hd__o22a_1
X_6984_ _1413_ _2691_ net357 _2692_ VGND VGND 
+ VPWR
+ VPWR _0262_ sky130_fd_sc_hd__o22a_1
X_6985_ \hkspi.wrstb\ \hkspi.rdstb\ _0079_ VGND VGND VPWR 
+ VPWR
+ _2693_ sky130_fd_sc_hd__o21ai_4
X_6986_ _1081_ _2693_ _1801_ VGND VGND VPWR 
+ VPWR
+ _0034_ sky130_fd_sc_hd__o21ai_1
X_6987_ _1082_ _2693_ _2689_ VGND VGND VPWR 
+ VPWR
+ _0035_ sky130_fd_sc_hd__o21ai_1
X_6988_ _1083_ _2693_ _2685_ VGND VGND VPWR 
+ VPWR
+ _0036_ sky130_fd_sc_hd__o21ai_1
X_6989_ _1084_ _2693_ _2681_ VGND VGND VPWR 
+ VPWR
+ _0037_ sky130_fd_sc_hd__o21ai_1
X_6990_ \hkspi.pre_pass_thru_user\ _1834_ _1426_ \hkspi.state[1]\ VGND VGND 
+ VPWR
+ VPWR _0029_ sky130_fd_sc_hd__a31o_1
X_6991_ serial_xfer VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__inv_2
X_6992_ _1666_ _1733_ \xfer_state[0]\ _2694_ VGND VGND 
+ VPWR
+ VPWR _0038_ sky130_fd_sc_hd__a2bb2o_1
X_6993_ \xfer_state[1]\ net306 \xfer_state[1]\ _1672_ \xfer_state[2]\ VGND 
+ VGND
+ VPWR VPWR _0039_ sky130_fd_sc_hd__a221o_2
X_6994_ _1708_ \pad_count_2[4]\ VGND VGND VPWR VPWR 
+ _2695_
+ sky130_fd_sc_hd__or2_4
X_6995_ \pad_count_2[3]\ _1714_ _1726_ VGND VGND VPWR 
+ VPWR
+ _2696_ sky130_fd_sc_hd__or3_1
X_6996_ _2695_ _2696_ VGND VGND VPWR VPWR 
+ _2697_
+ sky130_fd_sc_hd__nor2_2
X_6997_ _1665_ net306 _1672_ VGND VGND VPWR 
+ VPWR
+ _2698_ sky130_fd_sc_hd__or3_2
X_6998_ _1688_ _2694_ _2697_ _2698_ VGND VGND 
+ VPWR
+ VPWR _0040_ sky130_fd_sc_hd__o22ai_2
X_6999__13 _2698_ VGND VGND VPWR VPWR net391 sky130_fd_sc_hd__inv_2
X_7000_ \xfer_state[3]\ _1733_ _2697_ net391 VGND VGND 
+ VPWR
+ VPWR _0041_ sky130_fd_sc_hd__a22o_2
X_7001_ \wbbd_state[6]\ _1799_ VGND VGND VPWR VPWR 
+ _2700_
+ sky130_fd_sc_hd__or2_1
X_7002_ _2700_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
X_7003_ _1423_ _1429_ _1138_ _0091_ VGND VGND 
+ VPWR
+ VPWR _2701_ sky130_fd_sc_hd__and4bb_1
X_7004_ _1127_ _1419_ _1820_ _0087_ _2701_ VGND 
+ VGND
+ VPWR VPWR _2702_ sky130_fd_sc_hd__o32a_1
X_7005_ _2702_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__inv_2
X_7006_ \hkspi.pre_pass_thru_mgmt\ _1420_ \hkspi.state[0]\ \hkspi.state[4]\ VGND VGND 
+ VPWR
+ VPWR _0032_ sky130_fd_sc_hd__a31o_1
X_7007_ _1425_ _1426_ _1834_ \hkspi.state[3]\ _1419_ VGND 
+ VGND
+ VPWR VPWR _0031_ sky130_fd_sc_hd__a32o_1
X_7008_ _1419_ _1820_ VGND VGND VPWR VPWR 
+ _2703_
+ sky130_fd_sc_hd__or2_1
X_7009_ \hkspi.state[3]\ _1420_ \hkspi.state[2]\ _2703_ VGND VGND 
+ VPWR
+ VPWR _0030_ sky130_fd_sc_hd__a22o_1
X_7010_ \hkspi.pass_thru_mgmt_delay\ net75 VGND VGND VPWR VPWR 
+ net253
+ sky130_fd_sc_hd__nor2_1
X_7011_ \hkspi.pass_thru_mgmt\ net75 VGND VGND VPWR VPWR 
+ net251
+ sky130_fd_sc_hd__nor2_1
X_7012_ \hkspi.pass_thru_mgmt_delay\ net86 VGND VGND VPWR VPWR 
+ _2704_
+ sky130_fd_sc_hd__or2b_1
X_7013_ _2704_ VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__clkbuf_1
X_7014_ net255 VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__inv_2
X_7015_ \hkspi.pass_thru_mgmt\ net88 VGND VGND VPWR VPWR 
+ _2705_
+ sky130_fd_sc_hd__or2_1
X_7016_ _2705_ VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__clkbuf_1
X_7017_ net259 VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__inv_2
X_7018_ \hkspi.pass_thru_mgmt_delay\ net73 VGND VGND VPWR VPWR 
+ _2706_
+ sky130_fd_sc_hd__and2b_1
X_7019_ _2706_ VGND VGND VPWR VPWR net312 sky130_fd_sc_hd__buf_6
X_7020_ \hkspi.pass_thru_mgmt\ net74 VGND VGND VPWR VPWR 
+ _2707_
+ sky130_fd_sc_hd__and2b_1
X_7021_ _2707_ VGND VGND VPWR VPWR net313 sky130_fd_sc_hd__buf_4
X_7022_ net380 _1125_ VGND VGND VPWR VPWR 
+ _0098_
+ sky130_fd_sc_hd__nor2_2
X_7023_ \pad_count_2[3]\ \pad_count_2[2]\ VGND VGND VPWR VPWR 
+ _2708_
+ sky130_fd_sc_hd__or2_2
X_7024_ \pad_count_2[1]\ \pad_count_2[0]\ _2708_ _2695_ VGND VGND 
+ VPWR
+ VPWR _2709_ sky130_fd_sc_hd__or4_1
X_7025_ _2709_ VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__buf_8
X_7026_ \pad_count_2[5]\ \pad_count_2[4]\ VGND VGND VPWR VPWR 
+ _2711_
+ sky130_fd_sc_hd__or2_1
X_7027_ _2711_ VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__clkbuf_4
X_7028_ _1712_ _2708_ VGND VGND VPWR VPWR 
+ _2713_
+ sky130_fd_sc_hd__or2_1
X_7029_ _2712_ _2713_ VGND VGND VPWR VPWR 
+ _2714_
+ sky130_fd_sc_hd__or2_1
X_7030_ _2714_ VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__buf_8
X_7031_ _1727_ _2708_ VGND VGND VPWR VPWR 
+ _2716_
+ sky130_fd_sc_hd__or2_1
X_7032_ _2712_ _2716_ VGND VGND VPWR VPWR 
+ _2717_
+ sky130_fd_sc_hd__or2_1
X_7033_ _2717_ VGND VGND VPWR VPWR _2718_ sky130_fd_sc_hd__buf_8
X_7034_ _1726_ _2708_ VGND VGND VPWR VPWR 
+ _2719_
+ sky130_fd_sc_hd__or2_1
X_7035_ _2719_ _2712_ VGND VGND VPWR VPWR 
+ _2720_
+ sky130_fd_sc_hd__or2_1
X_7036_ _2720_ VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__buf_6
X_7037_ _1713_ \pad_count_2[2]\ VGND VGND VPWR VPWR 
+ _2722_
+ sky130_fd_sc_hd__or2_2
X_7038_ \pad_count_2[1]\ \pad_count_2[0]\ _2722_ _2712_ VGND VGND 
+ VPWR
+ VPWR _2723_ sky130_fd_sc_hd__or4_1
X_7039_ _2723_ VGND VGND VPWR VPWR _2724_ sky130_fd_sc_hd__clkbuf_16
X_7040_ _2715_ _2718_ _2721_ _2724_ VGND VGND 
+ VPWR
+ VPWR _2725_ sky130_fd_sc_hd__and4_1
X_7041_ _1716_ _2712_ VGND VGND VPWR VPWR 
+ _2726_
+ sky130_fd_sc_hd__or2_4
X_7042_ _1727_ _2722_ _2712_ VGND VGND VPWR 
+ VPWR
+ _2727_ sky130_fd_sc_hd__or3_1
X_7043_ _2727_ VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__buf_8
X_7044_ _2695_ _2719_ VGND VGND VPWR VPWR 
+ _2729_
+ sky130_fd_sc_hd__or2_1
X_7045_ _2729_ VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__buf_8
X_7046_ _1726_ _2722_ _2712_ VGND VGND VPWR 
+ VPWR
+ _2731_ sky130_fd_sc_hd__or3_1
X_7047_ _2731_ VGND VGND VPWR VPWR _2732_ sky130_fd_sc_hd__clkbuf_16
X_7048_ _2726_ _2728_ _2730_ _2732_ VGND VGND 
+ VPWR
+ VPWR _2733_ sky130_fd_sc_hd__and4_1
X_7049_ _1715_ _1726_ _2712_ VGND VGND VPWR 
+ VPWR
+ _2734_ sky130_fd_sc_hd__or3_1
X_7050_ _2734_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__buf_8
X_7051_ \pad_count_2[3]\ _1714_ _1727_ VGND VGND VPWR 
+ VPWR
+ _2736_ sky130_fd_sc_hd__or3_1
X_7052_ _2695_ _2736_ VGND VGND VPWR VPWR 
+ _2737_
+ sky130_fd_sc_hd__or2_1
X_7053_ _2737_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__buf_8
X_7054_ _2696_ _2712_ VGND VGND VPWR VPWR 
+ _2739_
+ sky130_fd_sc_hd__or2_1
X_7055_ _2739_ VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__buf_6
X_7056_ \pad_count_2[3]\ _1714_ \pad_count_2[1]\ \pad_count_2[0]\ VGND VGND 
+ VPWR
+ VPWR _2741_ sky130_fd_sc_hd__or4_1
X_7057_ _2712_ _2741_ VGND VGND VPWR VPWR 
+ _2742_
+ sky130_fd_sc_hd__or2_1
X_7058_ _2742_ VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__buf_8
X_7059_ _2735_ _2738_ _2740_ _2743_ VGND VGND 
+ VPWR
+ VPWR _2744_ sky130_fd_sc_hd__and4_1
X_7060_ _1712_ _2722_ _2712_ VGND VGND VPWR 
+ VPWR
+ _2745_ sky130_fd_sc_hd__or3_1
X_7061_ _2745_ VGND VGND VPWR VPWR _2746_ sky130_fd_sc_hd__buf_8
X_7062_ _2695_ _2741_ VGND VGND VPWR VPWR 
+ _2747_
+ sky130_fd_sc_hd__or2_1
X_7063_ _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__buf_8
X_7064_ _2695_ _2716_ VGND VGND VPWR VPWR 
+ _2749_
+ sky130_fd_sc_hd__or2_1
X_7065_ _2749_ VGND VGND VPWR VPWR _2750_ sky130_fd_sc_hd__buf_8
X_7066_ \pad_count_2[1]\ \pad_count_2[0]\ _1715_ _2712_ VGND VGND 
+ VPWR
+ VPWR _2751_ sky130_fd_sc_hd__or4_1
X_7067_ _2751_ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__clkbuf_16
X_7068_ _2746_ _2748_ _2750_ _2752_ VGND VGND 
+ VPWR
+ VPWR _2753_ sky130_fd_sc_hd__and4_1
X_7069_ _2712_ _2736_ VGND VGND VPWR VPWR 
+ _2754_
+ sky130_fd_sc_hd__or2_1
X_7070_ _2754_ VGND VGND VPWR VPWR _2755_ sky130_fd_sc_hd__buf_8
X_7071_ _1724_ _2712_ VGND VGND VPWR VPWR 
+ _2756_
+ sky130_fd_sc_hd__or2_1
X_7072_ _2756_ VGND VGND VPWR VPWR _2757_ sky130_fd_sc_hd__buf_8
X_7073_ _1715_ _1727_ _2712_ VGND VGND VPWR 
+ VPWR
+ _2758_ sky130_fd_sc_hd__or3_1
X_7074_ _2758_ VGND VGND VPWR VPWR _2759_ sky130_fd_sc_hd__buf_8
X_7075_ _2695_ _2713_ VGND VGND VPWR VPWR 
+ _2760_
+ sky130_fd_sc_hd__or2_1
X_7076_ _2760_ VGND VGND VPWR VPWR _2761_ sky130_fd_sc_hd__buf_8
X_7077_ _2755_ _2757_ _2759_ _2761_ VGND VGND 
+ VPWR
+ VPWR _2762_ sky130_fd_sc_hd__and4_1
X_7078_ _2733_ _2744_ _2753_ _2762_ VGND VGND 
+ VPWR
+ VPWR _2763_ sky130_fd_sc_hd__and4_1
X_7079_ _1719_ _2710_ _2725_ _2763_ VGND VGND 
+ VPWR
+ VPWR _2764_ sky130_fd_sc_hd__and4_1
X_7080_ _2764_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__buf_6
X_7081_ _1715_ _1727_ _1719_ VGND VGND VPWR 
+ VPWR
+ _2765_ sky130_fd_sc_hd__or3_1
X_7082_ _2765_ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__buf_8
X_7083_ _1715_ _1726_ _1719_ VGND VGND VPWR 
+ VPWR
+ _2767_ sky130_fd_sc_hd__or3_1
X_7084_ _2767_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__buf_8
X_7085_ _1719_ _2736_ VGND VGND VPWR VPWR 
+ _2769_
+ sky130_fd_sc_hd__or2_1
X_7086_ _2769_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__buf_8
X_7087_ _1719_ _2741_ VGND VGND VPWR VPWR 
+ _2771_
+ sky130_fd_sc_hd__or2_1
X_7088_ _2771_ VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__buf_8
X_7089_ _1393_ _2770_ _1391_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2773_ sky130_fd_sc_hd__o22a_1
X_7090_ _1199_ _2759_ _1230_ _2761_ _2773_ VGND 
+ VGND
+ VPWR VPWR _2774_ sky130_fd_sc_hd__o221a_1
X_7091_ _1333_ _2766_ _1328_ _2768_ _2774_ VGND 
+ VGND
+ VPWR VPWR _2775_ sky130_fd_sc_hd__o221a_1
X_7092_ _1252_ _2721_ _1143_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2776_ sky130_fd_sc_hd__o22a_1
X_7093_ _1219_ _2728_ _1180_ _2755_ _2776_ VGND 
+ VGND
+ VPWR VPWR _2777_ sky130_fd_sc_hd__o221a_1
X_7094_ _1719_ _2696_ VGND VGND VPWR VPWR 
+ _2778_
+ sky130_fd_sc_hd__or2_1
X_7095_ _2778_ VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__buf_8
X_7096_ _1719_ _1724_ VGND VGND VPWR VPWR 
+ _2780_
+ sky130_fd_sc_hd__or2_1
X_7097_ _2780_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__buf_8
X_7098_ \pad_count_2[1]\ \pad_count_2[0]\ _1715_ _1719_ VGND VGND 
+ VPWR
+ VPWR _2782_ sky130_fd_sc_hd__or4_1
X_7099_ _2782_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__buf_8
X_7100_ _1403_ _2781_ _1387_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2784_ sky130_fd_sc_hd__o22a_1
X_7101_ _1374_ _2779_ _1258_ _2752_ _2784_ VGND 
+ VGND
+ VPWR VPWR _2785_ sky130_fd_sc_hd__o221a_1
X_7102_ _1311_ _2710_ _1205_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2786_ sky130_fd_sc_hd__o22a_1
X_7103_ _1211_ _2738_ _1223_ _2750_ _2786_ VGND 
+ VGND
+ VPWR VPWR _2787_ sky130_fd_sc_hd__o221a_1
X_7104_ _1712_ _2722_ _1719_ VGND VGND VPWR 
+ VPWR
+ _2788_ sky130_fd_sc_hd__or3_1
X_7105_ _2788_ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__buf_8
X_7106_ _1187_ _2746_ _1272_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2790_ sky130_fd_sc_hd__o22a_1
X_7107_ _1213_ _2732_ _1248_ _2718_ _2790_ VGND 
+ VGND
+ VPWR VPWR _2791_ sky130_fd_sc_hd__o221a_1
X_7108_ _2777_ _2785_ _2787_ _2791_ VGND VGND 
+ VPWR
+ VPWR _2792_ sky130_fd_sc_hd__and4_1
X_7109_ _1719_ _2716_ VGND VGND VPWR VPWR 
+ _2793_
+ sky130_fd_sc_hd__or2_1
X_7110_ _2793_ VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__buf_8
X_7111_ \pad_count_2[1]\ \pad_count_2[0]\ _2708_ _1719_ VGND VGND 
+ VPWR
+ VPWR _2795_ sky130_fd_sc_hd__or4_2
X_7112_ _2795_ VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__buf_8
X_7113_ _1221_ _2796_ _1147_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2797_ sky130_fd_sc_hd__o22a_1
X_7114_ _1195_ _2724_ _1283_ _2794_ _2797_ VGND 
+ VGND
+ VPWR VPWR _2798_ sky130_fd_sc_hd__o221a_1
X_7115_ _1719_ _2719_ VGND VGND VPWR VPWR 
+ _2799_
+ sky130_fd_sc_hd__or2_1
X_7116_ _2799_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__buf_8
X_7117_ \pad_count_2[1]\ \pad_count_2[0]\ _2722_ _1719_ VGND VGND 
+ VPWR
+ VPWR _2801_ sky130_fd_sc_hd__or4_1
X_7118_ _2801_ VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__buf_8
X_7119_ _1324_ _2802_ _1154_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2803_ sky130_fd_sc_hd__o22a_1
X_7120_ _1166_ _2743_ _1354_ _2800_ _2803_ VGND 
+ VGND
+ VPWR VPWR _2804_ sky130_fd_sc_hd__o221a_1
X_7121_ _1238_ _2726_ VGND VGND VPWR VPWR 
+ _2805_
+ sky130_fd_sc_hd__or2_1
X_7122_ _1294_ _1721_ _1320_ _2715_ _2805_ VGND 
+ VGND
+ VPWR VPWR _2806_ sky130_fd_sc_hd__o221a_1
X_7123_ _1719_ _2713_ VGND VGND VPWR VPWR 
+ _2807_
+ sky130_fd_sc_hd__or2_1
X_7124_ _2807_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__buf_8
X_7125_ _1726_ _2722_ _1719_ VGND VGND VPWR 
+ VPWR
+ _2809_ sky130_fd_sc_hd__or3_1
X_7126_ _2809_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__buf_8
X_7127_ _1727_ _2722_ _1719_ VGND VGND VPWR 
+ VPWR
+ _2811_ sky130_fd_sc_hd__or3_1
X_7128_ _2811_ VGND VGND VPWR VPWR _2812_ sky130_fd_sc_hd__buf_8
X_7129_ _1292_ _2810_ _1335_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2813_ sky130_fd_sc_hd__o22a_1
X_7130_ _1405_ _2808_ _1250_ _2748_ _2813_ VGND 
+ VGND
+ VPWR VPWR _2814_ sky130_fd_sc_hd__o221a_1
X_7131_ _2798_ _2804_ _2806_ _2814_ VGND VGND 
+ VPWR
+ VPWR _2815_ sky130_fd_sc_hd__and4_1
X_7132_ _2775_ _2792_ _2815_ VGND VGND VPWR 
+ VPWR
+ _2816_ sky130_fd_sc_hd__and3_4
X_7133_ _2816_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_7134_ _2588_ _2770_ _2590_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2817_ sky130_fd_sc_hd__o22a_1
X_7135_ _2626_ _2759_ _2651_ _2761_ _2817_ VGND 
+ VGND
+ VPWR VPWR _2818_ sky130_fd_sc_hd__o221a_1
X_7136_ _2560_ _2766_ _2522_ _2768_ _2818_ VGND 
+ VGND
+ VPWR VPWR _2819_ sky130_fd_sc_hd__o221a_1
X_7137_ _2645_ _2721_ _2534_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2820_ sky130_fd_sc_hd__o22a_1
X_7138_ _2668_ _2728_ _2656_ _2755_ _2820_ VGND 
+ VGND
+ VPWR VPWR _2821_ sky130_fd_sc_hd__o221a_1
X_7139_ _2589_ _2781_ _2567_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2822_ sky130_fd_sc_hd__o22a_1
X_7140_ _2600_ _2779_ _2674_ _2752_ _2822_ VGND 
+ VGND
+ VPWR VPWR _2823_ sky130_fd_sc_hd__o221a_1
X_7141_ _2554_ _2710_ _2661_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2824_ sky130_fd_sc_hd__o22a_1
X_7142_ _2649_ _2738_ _2640_ _2750_ _2824_ VGND 
+ VGND
+ VPWR VPWR _2825_ sky130_fd_sc_hd__o221a_1
X_7143_ _2625_ _2746_ _2595_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2826_ sky130_fd_sc_hd__o22a_1
X_7144_ _2614_ _2732_ _2643_ _2718_ _2826_ VGND 
+ VGND
+ VPWR VPWR _2827_ sky130_fd_sc_hd__o221a_1
X_7145_ _2821_ _2823_ _2825_ _2827_ VGND VGND 
+ VPWR
+ VPWR _2828_ sky130_fd_sc_hd__and4_1
X_7146_ _2630_ _2796_ _2624_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2829_ sky130_fd_sc_hd__o22a_1
X_7147_ _2655_ _2724_ _2528_ _2794_ _2829_ VGND 
+ VGND
+ VPWR VPWR _2830_ sky130_fd_sc_hd__o221a_1
X_7148_ _2523_ _2802_ _2650_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2831_ sky130_fd_sc_hd__o22a_1
X_7149_ _2654_ _2743_ _2594_ _2800_ _2831_ VGND 
+ VGND
+ VPWR VPWR _2832_ sky130_fd_sc_hd__o221a_1
X_7150_ _2615_ _2726_ VGND VGND VPWR VPWR 
+ _2833_
+ sky130_fd_sc_hd__or2_1
X_7151_ _2553_ _1721_ _2648_ _2715_ _2833_ VGND 
+ VGND
+ VPWR VPWR _2834_ sky130_fd_sc_hd__o221a_1
X_7152_ _2558_ _2810_ _2579_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2835_ sky130_fd_sc_hd__o22a_1
X_7153_ _2606_ _2808_ _2619_ _2748_ _2835_ VGND 
+ VGND
+ VPWR VPWR _2836_ sky130_fd_sc_hd__o221a_1
X_7154_ _2830_ _2832_ _2834_ _2836_ VGND VGND 
+ VPWR
+ VPWR _2837_ sky130_fd_sc_hd__and4_1
X_7155_ _2819_ _2828_ _2837_ VGND VGND VPWR 
+ VPWR
+ _0103_ sky130_fd_sc_hd__nand3_4
X_7156_ _2450_ _2770_ _2447_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2838_ sky130_fd_sc_hd__o22a_1
X_7157_ _2401_ _2759_ _2430_ _2761_ _2838_ VGND 
+ VGND
+ VPWR VPWR _2839_ sky130_fd_sc_hd__o221a_1
X_7158_ _2454_ _2766_ _2441_ _2768_ _2839_ VGND 
+ VGND
+ VPWR VPWR _2840_ sky130_fd_sc_hd__o221a_1
X_7159_ _2404_ _2721_ _2491_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2841_ sky130_fd_sc_hd__o22a_1
X_7160_ _2381_ _2728_ _2418_ _2755_ _2841_ VGND 
+ VGND
+ VPWR VPWR _2842_ sky130_fd_sc_hd__o221a_1
X_7161_ _2497_ _2781_ _2472_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2843_ sky130_fd_sc_hd__o22a_1
X_7162_ _2473_ _2779_ _2380_ _2752_ _2843_ VGND 
+ VGND
+ VPWR VPWR _2844_ sky130_fd_sc_hd__o221a_1
X_7163_ _2457_ _2710_ _2370_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2845_ sky130_fd_sc_hd__o22a_1
X_7164_ _2485_ _2738_ _2490_ _2750_ _2845_ VGND 
+ VGND
+ VPWR VPWR _2846_ sky130_fd_sc_hd__o221a_1
X_7165_ _2376_ _2746_ _2498_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2847_ sky130_fd_sc_hd__o22a_1
X_7166_ _2374_ _2732_ _2510_ _2718_ _2847_ VGND 
+ VGND
+ VPWR VPWR _2848_ sky130_fd_sc_hd__o221a_1
X_7167_ _2842_ _2844_ _2846_ _2848_ VGND VGND 
+ VPWR
+ VPWR _2849_ sky130_fd_sc_hd__and4_1
X_7168_ _2398_ _2796_ _2492_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2850_ sky130_fd_sc_hd__o22a_1
X_7169_ _2424_ _2724_ _2474_ _2794_ _2850_ VGND 
+ VGND
+ VPWR VPWR _2851_ sky130_fd_sc_hd__o221a_1
X_7170_ _2431_ _2802_ _2423_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2852_ sky130_fd_sc_hd__o22a_1
X_7171_ _2512_ _2743_ _2461_ _2800_ _2852_ VGND 
+ VGND
+ VPWR VPWR _2853_ sky130_fd_sc_hd__o221a_1
X_7172_ _2368_ _2726_ VGND VGND VPWR VPWR 
+ _2854_
+ sky130_fd_sc_hd__or2_1
X_7173_ _2500_ _1721_ _2410_ _2715_ _2854_ VGND 
+ VGND
+ VPWR VPWR _2855_ sky130_fd_sc_hd__o221a_1
X_7174_ _2387_ _2810_ _2429_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2856_ sky130_fd_sc_hd__o22a_1
X_7175_ _2504_ _2808_ _2475_ _2748_ _2856_ VGND 
+ VGND
+ VPWR VPWR _2857_ sky130_fd_sc_hd__o221a_1
X_7176_ _2851_ _2853_ _2855_ _2857_ VGND VGND 
+ VPWR
+ VPWR _2858_ sky130_fd_sc_hd__and4_1
X_7177_ _2840_ _2849_ _2858_ VGND VGND VPWR 
+ VPWR
+ _0105_ sky130_fd_sc_hd__nand3_4
X_7178_ _4427_ _2770_ _4426_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2859_ sky130_fd_sc_hd__o22a_1
X_7179_ _4419_ _2759_ _0094_ _2761_ _2859_ VGND 
+ VGND
+ VPWR VPWR _2860_ sky130_fd_sc_hd__o221a_1
X_7180_ _4435_ _2766_ _4436_ _2768_ _2860_ VGND 
+ VGND
+ VPWR VPWR _2861_ sky130_fd_sc_hd__o221a_2
X_7181_ _4408_ _2721_ _4412_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2862_ sky130_fd_sc_hd__o22a_1
X_7182_ _4415_ _2728_ _4411_ _2755_ _2862_ VGND 
+ VGND
+ VPWR VPWR _2863_ sky130_fd_sc_hd__o221a_1
X_7183_ _4429_ _2781_ _4434_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2864_ sky130_fd_sc_hd__o22a_1
X_7184_ _4428_ _2779_ _4418_ _2752_ _2864_ VGND 
+ VGND
+ VPWR VPWR _2865_ sky130_fd_sc_hd__o221a_1
X_7185_ _4438_ _2710_ _4420_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2866_ sky130_fd_sc_hd__o22a_1
X_7186_ _0092_ _2738_ _4439_ _2750_ _2866_ VGND 
+ VGND
+ VPWR VPWR _2867_ sky130_fd_sc_hd__o221a_2
X_7187_ _4417_ _2746_ _4433_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2868_ sky130_fd_sc_hd__o22a_1
X_7188_ _4416_ _2732_ _2280_ _2718_ _2868_ VGND 
+ VGND
+ VPWR VPWR _2869_ sky130_fd_sc_hd__o221a_1
X_7189_ _2863_ _2865_ _2867_ _2869_ VGND VGND 
+ VPWR
+ VPWR _2870_ sky130_fd_sc_hd__and4_1
X_7190_ _4422_ _2796_ _4413_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2871_ sky130_fd_sc_hd__o22a_1
X_7191_ _4414_ _2724_ _4423_ _2794_ _2871_ VGND 
+ VGND
+ VPWR VPWR _2872_ sky130_fd_sc_hd__o221a_1
X_7192_ _4430_ _2802_ _4440_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2873_ sky130_fd_sc_hd__o22a_1
X_7193_ _4410_ _2743_ _4424_ _2800_ _2873_ VGND 
+ VGND
+ VPWR VPWR _2874_ sky130_fd_sc_hd__o221a_1
X_7194_ _4421_ _2726_ VGND VGND VPWR VPWR 
+ _2875_
+ sky130_fd_sc_hd__or2_1
X_7195_ _4437_ _1721_ _4409_ _2715_ _2875_ VGND 
+ VGND
+ VPWR VPWR _2876_ sky130_fd_sc_hd__o221a_1
X_7196_ _4432_ _2810_ _4431_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2877_ sky130_fd_sc_hd__o22a_1
X_7197_ _4425_ _2808_ _0093_ _2748_ _2877_ VGND 
+ VGND
+ VPWR VPWR _2878_ sky130_fd_sc_hd__o221a_1
X_7198_ _2872_ _2874_ _2876_ _2878_ VGND VGND 
+ VPWR
+ VPWR _2879_ sky130_fd_sc_hd__and4_1
X_7199_ _2861_ _2870_ _2879_ VGND VGND VPWR 
+ VPWR
+ _0107_ sky130_fd_sc_hd__nand3_4
X_7200_ _2193_ _2770_ _2135_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2880_ sky130_fd_sc_hd__o22a_1
X_7201_ _2149_ _2759_ _2239_ _2761_ _2880_ VGND 
+ VGND
+ VPWR VPWR _2881_ sky130_fd_sc_hd__o221a_1
X_7202_ _2205_ _2766_ _2168_ _2768_ _2881_ VGND 
+ VGND
+ VPWR VPWR _2882_ sky130_fd_sc_hd__o221a_2
X_7203_ _2241_ _2721_ _2115_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2883_ sky130_fd_sc_hd__o22a_1
X_7204_ _2131_ _2728_ _2240_ _2755_ _2883_ VGND 
+ VGND
+ VPWR VPWR _2884_ sky130_fd_sc_hd__o221a_1
X_7205_ _2107_ _2781_ _2127_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2885_ sky130_fd_sc_hd__o22a_1
X_7206_ _2174_ _2779_ _2146_ _2752_ _2885_ VGND 
+ VGND
+ VPWR VPWR _2886_ sky130_fd_sc_hd__o221a_1
X_7207_ _2206_ _2710_ _2155_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2887_ sky130_fd_sc_hd__o22a_1
X_7208_ _2134_ _2738_ _2170_ _2750_ _2887_ VGND 
+ VGND
+ VPWR VPWR _2888_ sky130_fd_sc_hd__o221a_1
X_7209_ _2150_ _2746_ _2180_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2889_ sky130_fd_sc_hd__o22a_1
X_7210_ _2145_ _2732_ _2217_ _2718_ _2889_ VGND 
+ VGND
+ VPWR VPWR _2890_ sky130_fd_sc_hd__o221a_1
X_7211_ _2884_ _2886_ _2888_ _2890_ VGND VGND 
+ VPWR
+ VPWR _2891_ sky130_fd_sc_hd__and4_1
X_7212_ _2138_ _2796_ _2246_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2892_ sky130_fd_sc_hd__o22a_1
X_7213_ _2235_ _2724_ _2176_ _2794_ _2892_ VGND 
+ VGND
+ VPWR VPWR _2893_ sky130_fd_sc_hd__o221a_1
X_7214_ _2124_ _2802_ _2214_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2894_ sky130_fd_sc_hd__o22a_1
X_7215_ _2234_ _2743_ _2199_ _2800_ _2894_ VGND 
+ VGND
+ VPWR VPWR _2895_ sky130_fd_sc_hd__o221a_1
X_7216_ _2158_ _2726_ VGND VGND VPWR VPWR 
+ _2896_
+ sky130_fd_sc_hd__or2_1
X_7217_ _2200_ _1721_ _2112_ _2715_ _2896_ VGND 
+ VGND
+ VPWR VPWR _2897_ sky130_fd_sc_hd__o221a_1
X_7218_ _2208_ _2810_ _2181_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2898_ sky130_fd_sc_hd__o22a_1
X_7219_ _2106_ _2808_ _2188_ _2748_ _2898_ VGND 
+ VGND
+ VPWR VPWR _2899_ sky130_fd_sc_hd__o221a_1
X_7220_ _2893_ _2895_ _2897_ _2899_ VGND VGND 
+ VPWR
+ VPWR _2900_ sky130_fd_sc_hd__and4_1
X_7221_ _2882_ _2891_ _2900_ VGND VGND VPWR 
+ VPWR
+ _0109_ sky130_fd_sc_hd__nand3_4
X_7222_ _2055_ _2770_ _2020_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2901_ sky130_fd_sc_hd__o22a_1
X_7223_ _2090_ _2759_ _2068_ _2761_ _2901_ VGND 
+ VGND
+ VPWR VPWR _2902_ sky130_fd_sc_hd__o221a_1
X_7224_ _2025_ _2766_ _2037_ _2768_ _2902_ VGND 
+ VGND
+ VPWR VPWR _2903_ sky130_fd_sc_hd__o221a_1
X_7225_ _2063_ _2721_ _2085_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2904_ sky130_fd_sc_hd__o22a_1
X_7226_ _2079_ _2728_ _2078_ _2755_ _2904_ VGND 
+ VGND
+ VPWR VPWR _2905_ sky130_fd_sc_hd__o221a_1
X_7227_ _2021_ _2781_ _2052_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2906_ sky130_fd_sc_hd__o22a_1
X_7228_ _2071_ _2779_ _2089_ _2752_ _2906_ VGND 
+ VGND
+ VPWR VPWR _2907_ sky130_fd_sc_hd__o221a_1
X_7229_ _2045_ _2710_ _2097_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2908_ sky130_fd_sc_hd__o22a_1
X_7230_ _2077_ _2738_ _2091_ _2750_ _2908_ VGND 
+ VGND
+ VPWR VPWR _2909_ sky130_fd_sc_hd__o221a_1
X_7231_ _2082_ _2746_ _2044_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2910_ sky130_fd_sc_hd__o22a_1
X_7232_ _2069_ _2732_ _2095_ _2718_ _2910_ VGND 
+ VGND
+ VPWR VPWR _2911_ sky130_fd_sc_hd__o221a_1
X_7233_ _2905_ _2907_ _2909_ _2911_ VGND VGND 
+ VPWR
+ VPWR _2912_ sky130_fd_sc_hd__and4_1
X_7234_ _2101_ _2796_ _2083_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2913_ sky130_fd_sc_hd__o22a_1
X_7235_ _2065_ _2724_ _2058_ _2794_ _2913_ VGND 
+ VGND
+ VPWR VPWR _2914_ sky130_fd_sc_hd__o221a_1
X_7236_ _2056_ _2802_ _2102_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2915_ sky130_fd_sc_hd__o22a_1
X_7237_ _2096_ _2743_ _2057_ _2800_ _2915_ VGND 
+ VGND
+ VPWR VPWR _2916_ sky130_fd_sc_hd__o221a_1
X_7238_ _2064_ _2726_ VGND VGND VPWR VPWR 
+ _2917_
+ sky130_fd_sc_hd__or2_1
X_7239_ _2027_ _1721_ _2084_ _2715_ _2917_ VGND 
+ VGND
+ VPWR VPWR _2918_ sky130_fd_sc_hd__o221a_1
X_7240_ _2072_ _2810_ _2022_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2919_ sky130_fd_sc_hd__o22a_1
X_7241_ _2050_ _2808_ _2092_ _2748_ _2919_ VGND 
+ VGND
+ VPWR VPWR _2920_ sky130_fd_sc_hd__o221a_1
X_7242_ _2914_ _2916_ _2918_ _2920_ VGND VGND 
+ VPWR
+ VPWR _2921_ sky130_fd_sc_hd__and4_1
X_7243_ _2903_ _2912_ _2921_ VGND VGND VPWR 
+ VPWR
+ _0111_ sky130_fd_sc_hd__nand3_4
X_7244_ _1943_ _2770_ _2008_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2922_ sky130_fd_sc_hd__o22a_1
X_7245_ _1961_ _2759_ _1935_ _2761_ _2922_ VGND 
+ VGND
+ VPWR VPWR _2923_ sky130_fd_sc_hd__o221a_1
X_7246_ _1944_ _2766_ _1978_ _2768_ _2923_ VGND 
+ VGND
+ VPWR VPWR _2924_ sky130_fd_sc_hd__o221a_1
X_7247_ _2015_ _2721_ _2007_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2925_ sky130_fd_sc_hd__o22a_1
X_7248_ _1958_ _2728_ _1998_ _2755_ _2925_ VGND 
+ VGND
+ VPWR VPWR _2926_ sky130_fd_sc_hd__o221a_1
X_7249_ _1952_ _2781_ _1951_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2927_ sky130_fd_sc_hd__o22a_1
X_7250_ _1979_ _2779_ _1966_ _2752_ _2927_ VGND 
+ VGND
+ VPWR VPWR _2928_ sky130_fd_sc_hd__o221a_1
X_7251_ _1973_ _2710_ _1962_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2929_ sky130_fd_sc_hd__o22a_1
X_7252_ _1953_ _2738_ _1984_ _2750_ _2929_ VGND 
+ VGND
+ VPWR VPWR _2930_ sky130_fd_sc_hd__o221a_1
X_7253_ _1965_ _2746_ _1982_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2931_ sky130_fd_sc_hd__o22a_1
X_7254_ _1967_ _2732_ _1941_ _2718_ _2931_ VGND 
+ VGND
+ VPWR VPWR _2932_ sky130_fd_sc_hd__o221a_1
X_7255_ _2926_ _2928_ _2930_ _2932_ VGND VGND 
+ VPWR
+ VPWR _2933_ sky130_fd_sc_hd__and4_1
X_7256_ _1959_ _2796_ _1995_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2934_ sky130_fd_sc_hd__o22a_1
X_7257_ _1977_ _2724_ _1938_ _2794_ _2934_ VGND 
+ VGND
+ VPWR VPWR _2935_ sky130_fd_sc_hd__o221a_1
X_7258_ _1954_ _2802_ _1988_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2936_ sky130_fd_sc_hd__o22a_1
X_7259_ _2001_ _2743_ _1936_ _2800_ _2936_ VGND 
+ VGND
+ VPWR VPWR _2937_ sky130_fd_sc_hd__o221a_1
X_7260_ _1964_ _2726_ VGND VGND VPWR VPWR 
+ _2938_
+ sky130_fd_sc_hd__or2_1
X_7261_ _1983_ _1721_ _2013_ _2715_ _2938_ VGND 
+ VGND
+ VPWR VPWR _2939_ sky130_fd_sc_hd__o221a_1
X_7262_ _1971_ _2810_ _1972_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2940_ sky130_fd_sc_hd__o22a_1
X_7263_ _1948_ _2808_ _1947_ _2748_ _2940_ VGND 
+ VGND
+ VPWR VPWR _2941_ sky130_fd_sc_hd__o221a_1
X_7264_ _2935_ _2937_ _2939_ _2941_ VGND VGND 
+ VPWR
+ VPWR _2942_ sky130_fd_sc_hd__and4_1
X_7265_ _2924_ _2933_ _2942_ VGND VGND VPWR 
+ VPWR
+ _0113_ sky130_fd_sc_hd__nand3_4
X_7266_ _1901_ _2770_ _1862_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2943_ sky130_fd_sc_hd__o22a_1
X_7267_ _1925_ _2759_ _1921_ _2761_ _2943_ VGND 
+ VGND
+ VPWR VPWR _2944_ sky130_fd_sc_hd__o221a_1
X_7268_ _1861_ _2766_ _1902_ _2768_ _2944_ VGND 
+ VGND
+ VPWR VPWR _2945_ sky130_fd_sc_hd__o221a_1
X_7269_ _1917_ _2721_ _1911_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2946_ sky130_fd_sc_hd__o22a_1
X_7270_ _1926_ _2728_ _1908_ _2755_ _2946_ VGND 
+ VGND
+ VPWR VPWR _2947_ sky130_fd_sc_hd__o221a_1
X_7271_ _1898_ _2781_ _1867_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2948_ sky130_fd_sc_hd__o22a_1
X_7272_ _1866_ _2779_ _1910_ _2752_ _2948_ VGND 
+ VGND
+ VPWR VPWR _2949_ sky130_fd_sc_hd__o221a_1
X_7273_ _1891_ _2710_ _1854_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2950_ sky130_fd_sc_hd__o22a_1
X_7274_ _1855_ _2738_ _1868_ _2750_ _2950_ VGND 
+ VGND
+ VPWR VPWR _2951_ sky130_fd_sc_hd__o221a_1
X_7275_ _1914_ _2746_ _1871_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2952_ sky130_fd_sc_hd__o22a_1
X_7276_ _1909_ _2732_ _1850_ _2718_ _2952_ VGND 
+ VGND
+ VPWR VPWR _2953_ sky130_fd_sc_hd__o221a_1
X_7277_ _2947_ _2949_ _2951_ _2953_ VGND VGND 
+ VPWR
+ VPWR _2954_ sky130_fd_sc_hd__and4_1
X_7278_ _1927_ _2796_ _1916_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2955_ sky130_fd_sc_hd__o22a_1
X_7279_ _1853_ _2724_ _1886_ _2794_ _2955_ VGND 
+ VGND
+ VPWR VPWR _2956_ sky130_fd_sc_hd__o221a_1
X_7280_ _1897_ _2802_ _1856_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2957_ sky130_fd_sc_hd__o22a_1
X_7281_ _1915_ _2743_ _1879_ _2800_ _2957_ VGND 
+ VGND
+ VPWR VPWR _2958_ sky130_fd_sc_hd__o221a_1
X_7282_ _1924_ _2726_ VGND VGND VPWR VPWR 
+ _2959_
+ sky130_fd_sc_hd__or2_1
X_7283_ _1860_ _1721_ _1847_ _2715_ _2959_ VGND 
+ VGND
+ VPWR VPWR _2960_ sky130_fd_sc_hd__o221a_1
X_7284_ _1892_ _2810_ _1904_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2961_ sky130_fd_sc_hd__o22a_1
X_7285_ _1878_ _2808_ _1849_ _2748_ _2961_ VGND 
+ VGND
+ VPWR VPWR _2962_ sky130_fd_sc_hd__o221a_1
X_7286_ _2956_ _2958_ _2960_ _2962_ VGND VGND 
+ VPWR
+ VPWR _2963_ sky130_fd_sc_hd__and4_1
X_7287_ _2945_ _2954_ _2963_ VGND VGND VPWR 
+ VPWR
+ _0115_ sky130_fd_sc_hd__nand3_4
X_7288_ _1376_ _2770_ _1326_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2964_ sky130_fd_sc_hd__o22a_1
X_7289_ _1207_ _2759_ _1150_ _2761_ _2964_ VGND 
+ VGND
+ VPWR VPWR _2965_ sky130_fd_sc_hd__o221a_1
X_7290_ _1365_ _2766_ _1343_ _2768_ _2965_ VGND 
+ VGND
+ VPWR VPWR _2966_ sky130_fd_sc_hd__o221a_1
X_7291_ _1156_ _2721_ _1254_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2967_ sky130_fd_sc_hd__o22a_1
X_7292_ _1240_ _2728_ _1263_ _2755_ _2967_ VGND 
+ VGND
+ VPWR VPWR _2968_ sky130_fd_sc_hd__o221a_1
X_7293_ _1407_ _2781_ _1360_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2969_ sky130_fd_sc_hd__o22a_1
X_7294_ _1401_ _2779_ _1201_ _2752_ _2969_ VGND 
+ VGND
+ VPWR VPWR _2970_ sky130_fd_sc_hd__o221a_1
X_7295_ _1379_ _2710_ _1185_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2971_ sky130_fd_sc_hd__o22a_1
X_7296_ _1228_ _2738_ _1367_ _2750_ _2971_ VGND 
+ VGND
+ VPWR VPWR _2972_ sky130_fd_sc_hd__o221a_2
X_7297_ _1191_ _2746_ _1314_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2973_ sky130_fd_sc_hd__o22a_1
X_7298_ _1164_ _2732_ _1301_ _2718_ _2973_ VGND 
+ VGND
+ VPWR VPWR _2974_ sky130_fd_sc_hd__o221a_1
X_7299_ _2968_ _2970_ _2972_ _2974_ VGND VGND 
+ VPWR
+ VPWR _2975_ sky130_fd_sc_hd__and4_1
X_7300_ _1197_ _2796_ _1178_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2976_ sky130_fd_sc_hd__o22a_1
X_7301_ _1173_ _2724_ _1139_ _2794_ _2976_ VGND 
+ VGND
+ VPWR VPWR _2977_ sky130_fd_sc_hd__o221a_2
X_7302_ _1279_ _2802_ _1265_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2978_ sky130_fd_sc_hd__o22a_1
X_7303_ _1244_ _2743_ _1397_ _2800_ _2978_ VGND 
+ VGND
+ VPWR VPWR _2979_ sky130_fd_sc_hd__o221a_1
X_7304_ _1189_ _2726_ VGND VGND VPWR VPWR 
+ _2980_
+ sky130_fd_sc_hd__or2_1
X_7305_ _1336_ _1721_ _1169_ _2715_ _2980_ VGND 
+ VGND
+ VPWR VPWR _2981_ sky130_fd_sc_hd__o221a_2
X_7306_ _1359_ _2810_ _1287_ _2812_ VGND VGND 
+ VPWR
+ VPWR _2982_ sky130_fd_sc_hd__o22a_1
X_7307_ _1395_ _2808_ _1242_ _2748_ _2982_ VGND 
+ VGND
+ VPWR VPWR _2983_ sky130_fd_sc_hd__o221a_1
X_7308_ _2977_ _2979_ _2981_ _2983_ VGND VGND 
+ VPWR
+ VPWR _2984_ sky130_fd_sc_hd__and4_1
X_7309_ _2966_ _2975_ _2984_ VGND VGND VPWR 
+ VPWR
+ _0117_ sky130_fd_sc_hd__nand3_4
X_7310_ _2608_ _2770_ _2602_ _2772_ VGND VGND 
+ VPWR
+ VPWR _2985_ sky130_fd_sc_hd__o22a_1
X_7311_ _2662_ _2759_ _2639_ _2761_ _2985_ VGND 
+ VGND
+ VPWR VPWR _2986_ sky130_fd_sc_hd__o221a_1
X_7312_ _2583_ _2766_ _2559_ _2768_ _2986_ VGND 
+ VGND
+ VPWR VPWR _2987_ sky130_fd_sc_hd__o221a_1
X_7313_ _2675_ _2721_ _2657_ _2740_ VGND VGND 
+ VPWR
+ VPWR _2988_ sky130_fd_sc_hd__o22a_1
X_7314_ _2618_ _2728_ _2535_ _2755_ _2988_ VGND 
+ VGND
+ VPWR VPWR _2989_ sky130_fd_sc_hd__o221a_1
X_7315_ _2578_ _2781_ _2580_ _2783_ VGND VGND 
+ VPWR
+ VPWR _2990_ sky130_fd_sc_hd__o22a_1
X_7316_ _2601_ _2779_ _2670_ _2752_ _2990_ VGND 
+ VGND
+ VPWR VPWR _2991_ sky130_fd_sc_hd__o221a_1
X_7317_ _2561_ _2710_ _2663_ _2735_ VGND VGND 
+ VPWR
+ VPWR _2992_ sky130_fd_sc_hd__o22a_1
X_7318_ _2537_ _2738_ _2575_ _2750_ _2992_ VGND 
+ VGND
+ VPWR VPWR _2993_ sky130_fd_sc_hd__o221a_1
X_7319_ _2667_ _2746_ _2540_ _2789_ VGND VGND 
+ VPWR
+ VPWR _2994_ sky130_fd_sc_hd__o22a_1
X_7320_ _2632_ _2732_ _2568_ _2718_ _2994_ VGND 
+ VGND
+ VPWR VPWR _2995_ sky130_fd_sc_hd__o221a_1
X_7321_ _2989_ _2991_ _2993_ _2995_ VGND VGND 
+ VPWR
+ VPWR _2996_ sky130_fd_sc_hd__and4_1
X_7322_ _2673_ _2796_ _2631_ _2757_ VGND VGND 
+ VPWR
+ VPWR _2997_ sky130_fd_sc_hd__o22a_1
X_7323_ _2644_ _2724_ _2633_ _2794_ _2997_ VGND 
+ VGND
+ VPWR VPWR _2998_ sky130_fd_sc_hd__o221a_2
X_7324_ _2609_ _2802_ _2627_ _2730_ VGND VGND 
+ VPWR
+ VPWR _2999_ sky130_fd_sc_hd__o22a_1
X_7325_ _2664_ _2743_ _2536_ _2800_ _2999_ VGND 
+ VGND
+ VPWR VPWR _3000_ sky130_fd_sc_hd__o221a_1
X_7326_ _2669_ _2726_ VGND VGND VPWR VPWR 
+ _3001_
+ sky130_fd_sc_hd__or2_1
X_7327_ _2591_ _1721_ _2637_ _2715_ _3001_ VGND 
+ VGND
+ VPWR VPWR _3002_ sky130_fd_sc_hd__o221a_2
X_7328_ _2547_ _2810_ _2603_ _2812_ VGND VGND 
+ VPWR
+ VPWR _3003_ sky130_fd_sc_hd__o22a_1
X_7329_ _2607_ _2808_ _2620_ _2748_ _3003_ VGND 
+ VGND
+ VPWR VPWR _3004_ sky130_fd_sc_hd__o221a_1
X_7330_ _2998_ _3000_ _3002_ _3004_ VGND VGND 
+ VPWR
+ VPWR _3005_ sky130_fd_sc_hd__and4_1
X_7331_ _2987_ _2996_ _3005_ VGND VGND VPWR 
+ VPWR
+ _0119_ sky130_fd_sc_hd__nand3_4
X_7332_ _2460_ _2770_ _2432_ _2772_ VGND VGND 
+ VPWR
+ VPWR _3006_ sky130_fd_sc_hd__o22a_1
X_7333_ _2382_ _2759_ _2493_ _2761_ _3006_ VGND 
+ VGND
+ VPWR VPWR _3007_ sky130_fd_sc_hd__o221a_1
X_7334_ _2467_ _2766_ _2442_ _2768_ _3007_ VGND 
+ VGND
+ VPWR VPWR _3008_ sky130_fd_sc_hd__o221a_1
X_7335_ _2469_ _2721_ _2480_ _2740_ VGND VGND 
+ VPWR
+ VPWR _3009_ sky130_fd_sc_hd__o22a_1
X_7336_ _2419_ _2728_ _2509_ _2755_ _3009_ VGND 
+ VGND
+ VPWR VPWR _3010_ sky130_fd_sc_hd__o221a_2
X_7337_ _2517_ _2781_ _2448_ _2783_ VGND VGND 
+ VPWR
+ VPWR _3011_ sky130_fd_sc_hd__o22a_1
X_7338_ _2466_ _2779_ _2375_ _2752_ _3011_ VGND 
+ VGND
+ VPWR VPWR _3012_ sky130_fd_sc_hd__o221a_1
X_7339_ _2394_ _2710_ _2371_ _2735_ VGND VGND 
+ VPWR
+ VPWR _3013_ sky130_fd_sc_hd__o22a_1
X_7340_ _2444_ _2738_ _2456_ _2750_ _3013_ VGND 
+ VGND
+ VPWR VPWR _3014_ sky130_fd_sc_hd__o221a_1
X_7341_ _2377_ _2746_ _2462_ _2789_ VGND VGND 
+ VPWR
+ VPWR _3015_ sky130_fd_sc_hd__o22a_2
X_7342_ _2383_ _2732_ _2482_ _2718_ _3015_ VGND 
+ VGND
+ VPWR VPWR _3016_ sky130_fd_sc_hd__o221a_1
X_7343_ _3010_ _3012_ _3014_ _3016_ VGND VGND 
+ VPWR
+ VPWR _3017_ sky130_fd_sc_hd__and4_1
X_7344_ _2369_ _2796_ _2487_ _2757_ VGND VGND 
+ VPWR
+ VPWR _3018_ sky130_fd_sc_hd__o22a_1
X_7345_ _2411_ _2724_ _2399_ _2794_ _3018_ VGND 
+ VGND
+ VPWR VPWR _3019_ sky130_fd_sc_hd__o221a_1
X_7346_ _2516_ _2802_ _2405_ _2730_ VGND VGND 
+ VPWR
+ VPWR _3020_ sky130_fd_sc_hd__o22a_1
X_7347_ _2468_ _2743_ _2455_ _2800_ _3020_ VGND 
+ VGND
+ VPWR VPWR _3021_ sky130_fd_sc_hd__o221a_1
X_7348_ _2400_ _2726_ VGND VGND VPWR VPWR 
+ _3022_
+ sky130_fd_sc_hd__or2_1
X_7349_ _2449_ _1721_ _2422_ _2715_ _3022_ VGND 
+ VGND
+ VPWR VPWR _3023_ sky130_fd_sc_hd__o221a_1
X_7350_ _2389_ _2810_ _2499_ _2812_ VGND VGND 
+ VPWR
+ VPWR _3024_ sky130_fd_sc_hd__o22a_1
X_7351_ _2437_ _2808_ _2438_ _2748_ _3024_ VGND 
+ VGND
+ VPWR VPWR _3025_ sky130_fd_sc_hd__o221a_2
X_7352_ _3019_ _3021_ _3023_ _3025_ VGND VGND 
+ VPWR
+ VPWR _3026_ sky130_fd_sc_hd__and4_1
X_7353_ _3008_ _3017_ _3026_ VGND VGND VPWR 
+ VPWR
+ _0121_ sky130_fd_sc_hd__nand3_4
X_7354_ _2313_ _2770_ _2354_ _2772_ VGND VGND 
+ VPWR
+ VPWR _3027_ sky130_fd_sc_hd__o22a_1
X_7355_ _2265_ _2759_ _2332_ _2761_ _3027_ VGND 
+ VGND
+ VPWR VPWR _3028_ sky130_fd_sc_hd__o221a_1
X_7356_ _2327_ _2766_ _2357_ _2768_ _3028_ VGND 
+ VGND
+ VPWR VPWR _3029_ sky130_fd_sc_hd__o221a_1
X_7357_ _2292_ _2721_ _2254_ _2740_ VGND VGND 
+ VPWR
+ VPWR _3030_ sky130_fd_sc_hd__o22a_1
X_7358_ _2271_ _2728_ _2297_ _2755_ _3030_ VGND 
+ VGND
+ VPWR VPWR _3031_ sky130_fd_sc_hd__o221a_2
X_7359_ _2349_ _2781_ _2307_ _2783_ VGND VGND 
+ VPWR
+ VPWR _3032_ sky130_fd_sc_hd__o22a_1
X_7360_ _2337_ _2779_ _2253_ _2752_ _3032_ VGND 
+ VGND
+ VPWR VPWR _3033_ sky130_fd_sc_hd__o221a_1
X_7361_ _2328_ _2710_ _2276_ _2735_ VGND VGND 
+ VPWR
+ VPWR _3034_ sky130_fd_sc_hd__o22a_1
X_7362_ _2284_ _2738_ _2314_ _2750_ _3034_ VGND 
+ VGND
+ VPWR VPWR _3035_ sky130_fd_sc_hd__o221a_1
X_7363_ _2331_ _2746_ _2344_ _2789_ VGND VGND 
+ VPWR
+ VPWR _3036_ sky130_fd_sc_hd__o22a_1
X_7364_ _2266_ _2732_ _2308_ _2718_ _3036_ VGND 
+ VGND
+ VPWR VPWR _3037_ sky130_fd_sc_hd__o221a_1
X_7365_ _3031_ _3033_ _3035_ _3037_ VGND VGND 
+ VPWR
+ VPWR _3038_ sky130_fd_sc_hd__and4_1
X_7366_ _2258_ _2796_ _2288_ _2757_ VGND VGND 
+ VPWR
+ VPWR _3039_ sky130_fd_sc_hd__o22a_1
X_7367_ _2259_ _2724_ _2275_ _2794_ _3039_ VGND 
+ VGND
+ VPWR VPWR _3040_ sky130_fd_sc_hd__o221a_1
X_7368_ _2350_ _2802_ _2270_ _2730_ VGND VGND 
+ VPWR
+ VPWR _3041_ sky130_fd_sc_hd__o22a_1
X_7369_ _2279_ _2743_ _2312_ _2800_ _3041_ VGND 
+ VGND
+ VPWR VPWR _3042_ sky130_fd_sc_hd__o221a_1
X_7370_ _2264_ _2726_ VGND VGND VPWR VPWR 
+ _3043_
+ sky130_fd_sc_hd__or2_1
X_7371_ _2301_ _1721_ _2289_ _2715_ _3043_ VGND 
+ VGND
+ VPWR VPWR _3044_ sky130_fd_sc_hd__o221a_1
X_7372_ _2306_ _2810_ _2353_ _2812_ VGND VGND 
+ VPWR
+ VPWR _3045_ sky130_fd_sc_hd__o22a_1
X_7373_ _2336_ _2808_ _2255_ _2748_ _3045_ VGND 
+ VGND
+ VPWR VPWR _3046_ sky130_fd_sc_hd__o221a_1
X_7374_ _3040_ _3042_ _3044_ _3046_ VGND VGND 
+ VPWR
+ VPWR _3047_ sky130_fd_sc_hd__and4_1
X_7375_ _3029_ _3038_ _3047_ VGND VGND VPWR 
+ VPWR
+ _0123_ sky130_fd_sc_hd__nand3_4
X_7376_ _2126_ _2770_ _2187_ _2772_ VGND VGND 
+ VPWR
+ VPWR _3048_ sky130_fd_sc_hd__o22a_1
X_7377_ _2140_ _2759_ _2218_ _2761_ _3048_ VGND 
+ VGND
+ VPWR VPWR _3049_ sky130_fd_sc_hd__o221a_1
X_7378_ _2175_ _2766_ _2165_ _2768_ _3049_ VGND 
+ VGND
+ VPWR VPWR _3050_ sky130_fd_sc_hd__o221a_1
X_7379_ _2242_ _2721_ _2109_ _2740_ VGND VGND 
+ VPWR
+ VPWR _3051_ sky130_fd_sc_hd__o22a_1
X_7380_ _2245_ _2728_ _2194_ _2755_ _3051_ VGND 
+ VGND
+ VPWR VPWR _3052_ sky130_fd_sc_hd__o221a_1
X_7381_ _2125_ _2781_ _2118_ _2783_ VGND VGND 
+ VPWR
+ VPWR _3053_ sky130_fd_sc_hd__o22a_1
X_7382_ _2177_ _2779_ _2152_ _2752_ _3053_ VGND 
+ VGND
+ VPWR VPWR _3054_ sky130_fd_sc_hd__o221a_1
X_7383_ _2195_ _2710_ _2157_ _2735_ VGND VGND 
+ VPWR
+ VPWR _3055_ sky130_fd_sc_hd__o22a_1
X_7384_ _2171_ _2738_ _2201_ _2750_ _3055_ VGND 
+ VGND
+ VPWR VPWR _3056_ sky130_fd_sc_hd__o221a_1
X_7385_ _2151_ _2746_ _2190_ _2789_ VGND VGND 
+ VPWR
+ VPWR _3057_ sky130_fd_sc_hd__o22a_1
X_7386_ _2147_ _2732_ _2223_ _2718_ _3057_ VGND 
+ VGND
+ VPWR VPWR _3058_ sky130_fd_sc_hd__o221a_1
X_7387_ _3052_ _3054_ _3056_ _3058_ VGND VGND 
+ VPWR
+ VPWR _3059_ sky130_fd_sc_hd__and4_1
X_7388_ _2139_ _2796_ _2219_ _2757_ VGND VGND 
+ VPWR
+ VPWR _3060_ sky130_fd_sc_hd__o22a_1
X_7389_ _2212_ _2724_ _2141_ _2794_ _3060_ VGND 
+ VGND
+ VPWR VPWR _3061_ sky130_fd_sc_hd__o221a_1
X_7390_ _2108_ _2802_ _2113_ _2730_ VGND VGND 
+ VPWR
+ VPWR _3062_ sky130_fd_sc_hd__o22a_1
X_7391_ _2236_ _2743_ _2202_ _2800_ _3062_ VGND 
+ VGND
+ VPWR VPWR _3063_ sky130_fd_sc_hd__o221a_1
X_7392_ _2156_ _2726_ VGND VGND VPWR VPWR 
+ _3064_
+ sky130_fd_sc_hd__or2_1
X_7393_ _2169_ _1721_ _2196_ _2715_ _3064_ VGND 
+ VGND
+ VPWR VPWR _3065_ sky130_fd_sc_hd__o221a_1
X_7394_ _2207_ _2810_ _2119_ _2812_ VGND VGND 
+ VPWR
+ VPWR _3066_ sky130_fd_sc_hd__o22a_1
X_7395_ _2182_ _2808_ _2121_ _2748_ _3066_ VGND 
+ VGND
+ VPWR VPWR _3067_ sky130_fd_sc_hd__o221a_1
X_7396_ _3061_ _3063_ _3065_ _3067_ VGND VGND 
+ VPWR
+ VPWR _3068_ sky130_fd_sc_hd__and4_1
X_7397_ _3050_ _3059_ _3068_ VGND VGND VPWR 
+ VPWR
+ _0125_ sky130_fd_sc_hd__nand3_4
X_7398_ _1693_ _1692_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _0127_ sky130_fd_sc_hd__nor3_4
X_7399_ _1702_ \pad_count_1[0]\ _1693_ _1695_ VGND VGND 
+ VPWR
+ VPWR _3069_ sky130_fd_sc_hd__or4_1
X_7400_ _3069_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__buf_6
X_7401_ \pad_count_1[1]\ _1703_ VGND VGND VPWR VPWR 
+ _3071_
+ sky130_fd_sc_hd__or2_4
X_7402_ \pad_count_1[3]\ VGND VGND VPWR VPWR _3072_ sky130_fd_sc_hd__inv_2
X_7403_ _3072_ _1699_ VGND VGND VPWR VPWR 
+ _3073_
+ sky130_fd_sc_hd__or2_4
X_7404_ _3071_ _3073_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3074_ sky130_fd_sc_hd__or3_1
X_7405_ _3074_ VGND VGND VPWR VPWR _3075_ sky130_fd_sc_hd__buf_6
X_7406_ \pad_count_1[3]\ _1699_ VGND VGND VPWR VPWR 
+ _3076_
+ sky130_fd_sc_hd__or2_4
X_7407_ _1702_ \pad_count_1[0]\ _3076_ _1695_ VGND VGND 
+ VPWR
+ VPWR _3077_ sky130_fd_sc_hd__or4_1
X_7408_ _3077_ VGND VGND VPWR VPWR _3078_ sky130_fd_sc_hd__buf_6
X_7409_ _1693_ _1704_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3079_ sky130_fd_sc_hd__or3_1
X_7410_ _3079_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__buf_6
X_7411_ _1374_ _3078_ _1320_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3081_ sky130_fd_sc_hd__o22a_1
X_7412_ _1354_ _3070_ _1199_ _3075_ _3081_ VGND 
+ VGND
+ VPWR VPWR _3082_ sky130_fd_sc_hd__o221a_1
X_7413_ _3072_ \pad_count_1[2]\ VGND VGND VPWR VPWR 
+ _3083_
+ sky130_fd_sc_hd__or2_4
X_7414_ _3083_ _1704_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3084_ sky130_fd_sc_hd__or3_1
X_7415_ _3084_ VGND VGND VPWR VPWR _3085_ sky130_fd_sc_hd__buf_6
X_7416_ _3071_ _3076_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3086_ sky130_fd_sc_hd__or3_1
X_7417_ _3086_ VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__buf_6
X_7418_ _1702_ \pad_count_1[0]\ _1693_ \pad_count_1[4]\ VGND VGND 
+ VPWR
+ VPWR _3088_ sky130_fd_sc_hd__or4_1
X_7419_ _3088_ VGND VGND VPWR VPWR _3089_ sky130_fd_sc_hd__buf_6
X_7420_ _3083_ _3071_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3090_ sky130_fd_sc_hd__or3_1
X_7421_ _3090_ VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__buf_6
X_7422_ _1252_ _3089_ _1335_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3092_ sky130_fd_sc_hd__o22a_1
X_7423_ _1187_ _3085_ _1180_ _3087_ _3092_ VGND 
+ VGND
+ VPWR VPWR _3093_ sky130_fd_sc_hd__o221a_1
X_7424_ _1692_ _3076_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3094_ sky130_fd_sc_hd__or3_1
X_7425_ _3094_ VGND VGND VPWR VPWR _3095_ sky130_fd_sc_hd__buf_8
X_7426_ _1704_ _3073_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3096_ sky130_fd_sc_hd__or3_1
X_7427_ _3096_ VGND VGND VPWR VPWR _3097_ sky130_fd_sc_hd__buf_8
X_7428_ _1294_ _3097_ _1221_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3098_ sky130_fd_sc_hd__o22a_1
X_7429_ _1702_ \pad_count_1[0]\ _3076_ \pad_count_1[4]\ VGND VGND 
+ VPWR
+ VPWR _3099_ sky130_fd_sc_hd__or4_1
X_7430_ _3099_ VGND VGND VPWR VPWR _3100_ sky130_fd_sc_hd__buf_6
X_7431_ _3083_ _1704_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3101_ sky130_fd_sc_hd__or3_1
X_7432_ _3101_ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__buf_6
X_7433_ _1692_ _3083_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3103_ sky130_fd_sc_hd__or3_1
X_7434_ _3103_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__buf_6
X_7435_ _1704_ _3076_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3105_ sky130_fd_sc_hd__or3_1
X_7436_ _3105_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__buf_6
X_7437_ _1324_ _3104_ _1403_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3107_ sky130_fd_sc_hd__o22a_1
X_7438_ _1143_ _3100_ _1272_ _3102_ _3107_ VGND 
+ VGND
+ VPWR VPWR _3108_ sky130_fd_sc_hd__o221a_1
X_7439_ _1166_ _3095_ _3098_ _3108_ VGND VGND 
+ VPWR
+ VPWR _3109_ sky130_fd_sc_hd__o211a_1
X_7440_ _1692_ _3073_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3110_ sky130_fd_sc_hd__or3_1
X_7441_ _3110_ VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__buf_8
X_7442_ _1702_ \pad_count_1[0]\ _3073_ _1695_ VGND VGND 
+ VPWR
+ VPWR _3112_ sky130_fd_sc_hd__or4_1
X_7443_ _3112_ VGND VGND VPWR VPWR _3113_ sky130_fd_sc_hd__buf_8
X_7444_ _1692_ _3076_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3114_ sky130_fd_sc_hd__or3_1
X_7445_ _3114_ VGND VGND VPWR VPWR _3115_ sky130_fd_sc_hd__buf_8
X_7446_ _1693_ _1704_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3116_ sky130_fd_sc_hd__or3_1
X_7447_ _3116_ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__buf_8
X_7448_ _1391_ _3115_ _1405_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3118_ sky130_fd_sc_hd__o22a_1
X_7449_ _1258_ _3111_ _1328_ _3113_ _3118_ VGND 
+ VGND
+ VPWR VPWR _3119_ sky130_fd_sc_hd__o221a_1
X_7450_ _3083_ _3071_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3120_ sky130_fd_sc_hd__or3_1
X_7451_ _3120_ VGND VGND VPWR VPWR _3121_ sky130_fd_sc_hd__buf_8
X_7452_ _3071_ _3076_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3122_ sky130_fd_sc_hd__or3_1
X_7453_ _3122_ VGND VGND VPWR VPWR _3123_ sky130_fd_sc_hd__buf_8
X_7454_ _1693_ _3071_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3124_ sky130_fd_sc_hd__or3_1
X_7455_ _3124_ VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__buf_8
X_7456_ _1693_ _3071_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3126_ sky130_fd_sc_hd__or3_1
X_7457_ _3126_ VGND VGND VPWR VPWR _3127_ sky130_fd_sc_hd__buf_8
X_7458_ _1283_ _3125_ _1248_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3128_ sky130_fd_sc_hd__o22a_1
X_7459_ _1219_ _3121_ _1393_ _3123_ _3128_ VGND 
+ VGND
+ VPWR VPWR _3129_ sky130_fd_sc_hd__o221a_1
X_7460_ _1692_ _3083_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3130_ sky130_fd_sc_hd__or3_1
X_7461_ _3130_ VGND VGND VPWR VPWR _3131_ sky130_fd_sc_hd__buf_8
X_7462_ _1692_ _3073_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3132_ sky130_fd_sc_hd__or3_1
X_7463_ _3132_ VGND VGND VPWR VPWR _3133_ sky130_fd_sc_hd__buf_8
X_7464_ _1702_ \pad_count_1[0]\ _3083_ \pad_count_1[4]\ VGND VGND 
+ VPWR
+ VPWR _3134_ sky130_fd_sc_hd__or4_1
X_7465_ _3134_ VGND VGND VPWR VPWR _3135_ sky130_fd_sc_hd__buf_8
X_7466_ _3071_ _3073_ _1695_ VGND VGND VPWR 
+ VPWR
+ _3136_ sky130_fd_sc_hd__or3_1
X_7467_ _3136_ VGND VGND VPWR VPWR _3137_ sky130_fd_sc_hd__buf_8
X_7468_ _1213_ _3135_ _1333_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3138_ sky130_fd_sc_hd__o22a_1
X_7469_ _1195_ _3131_ _1387_ _3133_ _3138_ VGND 
+ VGND
+ VPWR VPWR _3139_ sky130_fd_sc_hd__o221a_1
X_7470_ _1704_ _3076_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3140_ sky130_fd_sc_hd__or3_1
X_7471_ _3140_ VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__buf_8
X_7472_ _1704_ _3073_ \pad_count_1[4]\ VGND VGND VPWR 
+ VPWR
+ _3142_ sky130_fd_sc_hd__or3_1
X_7473_ _3142_ VGND VGND VPWR VPWR _3143_ sky130_fd_sc_hd__buf_8
X_7474_ _1702_ \pad_count_1[0]\ _3083_ _1695_ VGND VGND 
+ VPWR
+ VPWR _3144_ sky130_fd_sc_hd__or4_1
X_7475_ _3144_ VGND VGND VPWR VPWR _3145_ sky130_fd_sc_hd__buf_8
X_7476_ _1702_ \pad_count_1[0]\ _3073_ \pad_count_1[4]\ VGND VGND 
+ VPWR
+ VPWR _3146_ sky130_fd_sc_hd__or4_1
X_7477_ _3146_ VGND VGND VPWR VPWR _3147_ sky130_fd_sc_hd__buf_6
X_7478_ _1292_ _3145_ _1205_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3148_ sky130_fd_sc_hd__o22a_1
X_7479_ _1147_ _3141_ _1238_ _3143_ _3148_ VGND 
+ VGND
+ VPWR VPWR _3149_ sky130_fd_sc_hd__o221a_1
X_7480_ _3119_ _3129_ _3139_ _3149_ VGND VGND 
+ VPWR
+ VPWR _3150_ sky130_fd_sc_hd__and4_1
X_7481_ _3082_ _3093_ _3109_ _3150_ VGND VGND 
+ VPWR
+ VPWR _3151_ sky130_fd_sc_hd__and4_2
X_7482_ _3151_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_7483_ _2600_ _3078_ _2648_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3152_ sky130_fd_sc_hd__o22a_1
X_7484_ _2594_ _3070_ _2626_ _3075_ _3152_ VGND 
+ VGND
+ VPWR VPWR _3153_ sky130_fd_sc_hd__o221a_1
X_7485_ _2645_ _3089_ _2579_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3154_ sky130_fd_sc_hd__o22a_1
X_7486_ _2625_ _3085_ _2656_ _3087_ _3154_ VGND 
+ VGND
+ VPWR VPWR _3155_ sky130_fd_sc_hd__o221a_1
X_7487_ _2553_ _3097_ _2630_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3156_ sky130_fd_sc_hd__o22a_1
X_7488_ _2523_ _3104_ _2589_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3157_ sky130_fd_sc_hd__o22a_1
X_7489_ _2534_ _3100_ _2595_ _3102_ _3157_ VGND 
+ VGND
+ VPWR VPWR _3158_ sky130_fd_sc_hd__o221a_1
X_7490_ _2654_ _3095_ _3156_ _3158_ VGND VGND 
+ VPWR
+ VPWR _3159_ sky130_fd_sc_hd__o211a_1
X_7491_ _2590_ _3115_ _2606_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3160_ sky130_fd_sc_hd__o22a_1
X_7492_ _2674_ _3111_ _2522_ _3113_ _3160_ VGND 
+ VGND
+ VPWR VPWR _3161_ sky130_fd_sc_hd__o221a_1
X_7493_ _2528_ _3125_ _2643_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3162_ sky130_fd_sc_hd__o22a_1
X_7494_ _2668_ _3121_ _2588_ _3123_ _3162_ VGND 
+ VGND
+ VPWR VPWR _3163_ sky130_fd_sc_hd__o221a_1
X_7495_ _2614_ _3135_ _2560_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3164_ sky130_fd_sc_hd__o22a_1
X_7496_ _2655_ _3131_ _2567_ _3133_ _3164_ VGND 
+ VGND
+ VPWR VPWR _3165_ sky130_fd_sc_hd__o221a_1
X_7497_ _2558_ _3145_ _2661_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3166_ sky130_fd_sc_hd__o22a_1
X_7498_ _2624_ _3141_ _2615_ _3143_ _3166_ VGND 
+ VGND
+ VPWR VPWR _3167_ sky130_fd_sc_hd__o221a_1
X_7499_ _3161_ _3163_ _3165_ _3167_ VGND VGND 
+ VPWR
+ VPWR _3168_ sky130_fd_sc_hd__and4_1
X_7500_ _3153_ _3155_ _3159_ _3168_ VGND VGND 
+ VPWR
+ VPWR _0130_ sky130_fd_sc_hd__nand4_4
X_7501_ _2473_ _3078_ _2410_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3169_ sky130_fd_sc_hd__o22a_1
X_7502_ _2461_ _3070_ _2401_ _3075_ _3169_ VGND 
+ VGND
+ VPWR VPWR _3170_ sky130_fd_sc_hd__o221a_1
X_7503_ _2404_ _3089_ _2429_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3171_ sky130_fd_sc_hd__o22a_1
X_7504_ _2376_ _3085_ _2418_ _3087_ _3171_ VGND 
+ VGND
+ VPWR VPWR _3172_ sky130_fd_sc_hd__o221a_1
X_7505_ _2500_ _3097_ _2398_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3173_ sky130_fd_sc_hd__o22a_1
X_7506_ _2431_ _3104_ _2497_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3174_ sky130_fd_sc_hd__o22a_1
X_7507_ _2491_ _3100_ _2498_ _3102_ _3174_ VGND 
+ VGND
+ VPWR VPWR _3175_ sky130_fd_sc_hd__o221a_1
X_7508_ _2512_ _3095_ _3173_ _3175_ VGND VGND 
+ VPWR
+ VPWR _3176_ sky130_fd_sc_hd__o211a_1
X_7509_ _2447_ _3115_ _2504_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3177_ sky130_fd_sc_hd__o22a_1
X_7510_ _2380_ _3111_ _2441_ _3113_ _3177_ VGND 
+ VGND
+ VPWR VPWR _3178_ sky130_fd_sc_hd__o221a_1
X_7511_ _2474_ _3125_ _2510_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3179_ sky130_fd_sc_hd__o22a_1
X_7512_ _2381_ _3121_ _2450_ _3123_ _3179_ VGND 
+ VGND
+ VPWR VPWR _3180_ sky130_fd_sc_hd__o221a_1
X_7513_ _2374_ _3135_ _2454_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3181_ sky130_fd_sc_hd__o22a_1
X_7514_ _2424_ _3131_ _2472_ _3133_ _3181_ VGND 
+ VGND
+ VPWR VPWR _3182_ sky130_fd_sc_hd__o221a_1
X_7515_ _2387_ _3145_ _2370_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3183_ sky130_fd_sc_hd__o22a_1
X_7516_ _2492_ _3141_ _2368_ _3143_ _3183_ VGND 
+ VGND
+ VPWR VPWR _3184_ sky130_fd_sc_hd__o221a_1
X_7517_ _3178_ _3180_ _3182_ _3184_ VGND VGND 
+ VPWR
+ VPWR _3185_ sky130_fd_sc_hd__and4_2
X_7518_ _3170_ _3172_ _3176_ _3185_ VGND VGND 
+ VPWR
+ VPWR _0132_ sky130_fd_sc_hd__nand4_4
X_7519_ _4424_ _3070_ _4419_ _3075_ VGND VGND 
+ VPWR
+ VPWR _3186_ sky130_fd_sc_hd__o22a_1
X_7520_ _4428_ _3078_ _4409_ _3080_ _3186_ VGND 
+ VGND
+ VPWR VPWR _3187_ sky130_fd_sc_hd__o221a_1
X_7521_ _4408_ _3089_ _4431_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3188_ sky130_fd_sc_hd__o22a_1
X_7522_ _4417_ _3085_ _4411_ _3087_ _3188_ VGND 
+ VGND
+ VPWR VPWR _3189_ sky130_fd_sc_hd__o221a_1
X_7523_ _4437_ _3097_ _4422_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3190_ sky130_fd_sc_hd__o22a_1
X_7524_ _4430_ _3104_ _4429_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3191_ sky130_fd_sc_hd__o22a_1
X_7525_ _4412_ _3100_ _4433_ _3102_ _3191_ VGND 
+ VGND
+ VPWR VPWR _3192_ sky130_fd_sc_hd__o221a_1
X_7526_ _4410_ _3095_ _3190_ _3192_ VGND VGND 
+ VPWR
+ VPWR _3193_ sky130_fd_sc_hd__o211a_1
X_7527_ _4426_ _3115_ _4425_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3194_ sky130_fd_sc_hd__o22a_1
X_7528_ _4418_ _3111_ _4436_ _3113_ _3194_ VGND 
+ VGND
+ VPWR VPWR _3195_ sky130_fd_sc_hd__o221a_1
X_7529_ _4423_ _3125_ _2280_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3196_ sky130_fd_sc_hd__o22a_1
X_7530_ _4415_ _3121_ _4427_ _3123_ _3196_ VGND 
+ VGND
+ VPWR VPWR _3197_ sky130_fd_sc_hd__o221a_1
X_7531_ _4416_ _3135_ _4435_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3198_ sky130_fd_sc_hd__o22a_1
X_7532_ _4414_ _3131_ _4434_ _3133_ _3198_ VGND 
+ VGND
+ VPWR VPWR _3199_ sky130_fd_sc_hd__o221a_1
X_7533_ _4432_ _3145_ _4420_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3200_ sky130_fd_sc_hd__o22a_1
X_7534_ _4413_ _3141_ _4421_ _3143_ _3200_ VGND 
+ VGND
+ VPWR VPWR _3201_ sky130_fd_sc_hd__o221a_1
X_7535_ _3195_ _3197_ _3199_ _3201_ VGND VGND 
+ VPWR
+ VPWR _3202_ sky130_fd_sc_hd__and4_1
X_7536_ _3187_ _3189_ _3193_ _3202_ VGND VGND 
+ VPWR
+ VPWR _0134_ sky130_fd_sc_hd__nand4_4
X_7537_ _2174_ _3078_ _2112_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3203_ sky130_fd_sc_hd__o22a_1
X_7538_ _2199_ _3070_ _2149_ _3075_ _3203_ VGND 
+ VGND
+ VPWR VPWR _3204_ sky130_fd_sc_hd__o221a_1
X_7539_ _2241_ _3089_ _2181_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3205_ sky130_fd_sc_hd__o22a_1
X_7540_ _2150_ _3085_ _2240_ _3087_ _3205_ VGND 
+ VGND
+ VPWR VPWR _3206_ sky130_fd_sc_hd__o221a_1
X_7541_ _2200_ _3097_ _2138_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3207_ sky130_fd_sc_hd__o22a_1
X_7542_ _2124_ _3104_ _2107_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3208_ sky130_fd_sc_hd__o22a_1
X_7543_ _2115_ _3100_ _2180_ _3102_ _3208_ VGND 
+ VGND
+ VPWR VPWR _3209_ sky130_fd_sc_hd__o221a_1
X_7544_ _2234_ _3095_ _3207_ _3209_ VGND VGND 
+ VPWR
+ VPWR _3210_ sky130_fd_sc_hd__o211a_1
X_7545_ _2135_ _3115_ _2106_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3211_ sky130_fd_sc_hd__o22a_1
X_7546_ _2146_ _3111_ _2168_ _3113_ _3211_ VGND 
+ VGND
+ VPWR VPWR _3212_ sky130_fd_sc_hd__o221a_1
X_7547_ _2176_ _3125_ _2217_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3213_ sky130_fd_sc_hd__o22a_1
X_7548_ _2131_ _3121_ _2193_ _3123_ _3213_ VGND 
+ VGND
+ VPWR VPWR _3214_ sky130_fd_sc_hd__o221a_1
X_7549_ _2145_ _3135_ _2205_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3215_ sky130_fd_sc_hd__o22a_1
X_7550_ _2235_ _3131_ _2127_ _3133_ _3215_ VGND 
+ VGND
+ VPWR VPWR _3216_ sky130_fd_sc_hd__o221a_1
X_7551_ _2208_ _3145_ _2155_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3217_ sky130_fd_sc_hd__o22a_1
X_7552_ _2246_ _3141_ _2158_ _3143_ _3217_ VGND 
+ VGND
+ VPWR VPWR _3218_ sky130_fd_sc_hd__o221a_1
X_7553_ _3212_ _3214_ _3216_ _3218_ VGND VGND 
+ VPWR
+ VPWR _3219_ sky130_fd_sc_hd__and4_1
X_7554_ _3204_ _3206_ _3210_ _3219_ VGND VGND 
+ VPWR
+ VPWR _0136_ sky130_fd_sc_hd__nand4_4
X_7555_ _2071_ _3078_ _2084_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3220_ sky130_fd_sc_hd__o22a_1
X_7556_ _2057_ _3070_ _2090_ _3075_ _3220_ VGND 
+ VGND
+ VPWR VPWR _3221_ sky130_fd_sc_hd__o221a_1
X_7557_ _2063_ _3089_ _2022_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3222_ sky130_fd_sc_hd__o22a_1
X_7558_ _2082_ _3085_ _2078_ _3087_ _3222_ VGND 
+ VGND
+ VPWR VPWR _3223_ sky130_fd_sc_hd__o221a_1
X_7559_ _2027_ _3097_ _2101_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3224_ sky130_fd_sc_hd__o22a_1
X_7560_ _2056_ _3104_ _2021_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3225_ sky130_fd_sc_hd__o22a_1
X_7561_ _2085_ _3100_ _2044_ _3102_ _3225_ VGND 
+ VGND
+ VPWR VPWR _3226_ sky130_fd_sc_hd__o221a_1
X_7562_ _2096_ _3095_ _3224_ _3226_ VGND VGND 
+ VPWR
+ VPWR _3227_ sky130_fd_sc_hd__o211a_1
X_7563_ _2020_ _3115_ _2050_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3228_ sky130_fd_sc_hd__o22a_1
X_7564_ _2089_ _3111_ _2037_ _3113_ _3228_ VGND 
+ VGND
+ VPWR VPWR _3229_ sky130_fd_sc_hd__o221a_1
X_7565_ _2058_ _3125_ _2095_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3230_ sky130_fd_sc_hd__o22a_1
X_7566_ _2079_ _3121_ _2055_ _3123_ _3230_ VGND 
+ VGND
+ VPWR VPWR _3231_ sky130_fd_sc_hd__o221a_1
X_7567_ _2069_ _3135_ _2025_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3232_ sky130_fd_sc_hd__o22a_1
X_7568_ _2065_ _3131_ _2052_ _3133_ _3232_ VGND 
+ VGND
+ VPWR VPWR _3233_ sky130_fd_sc_hd__o221a_1
X_7569_ _2072_ _3145_ _2097_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3234_ sky130_fd_sc_hd__o22a_1
X_7570_ _2083_ _3141_ _2064_ _3143_ _3234_ VGND 
+ VGND
+ VPWR VPWR _3235_ sky130_fd_sc_hd__o221a_1
X_7571_ _3229_ _3231_ _3233_ _3235_ VGND VGND 
+ VPWR
+ VPWR _3236_ sky130_fd_sc_hd__and4_2
X_7572_ _3221_ _3223_ _3227_ _3236_ VGND VGND 
+ VPWR
+ VPWR _0138_ sky130_fd_sc_hd__nand4_4
X_7573_ _1979_ _3078_ _2013_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3237_ sky130_fd_sc_hd__o22a_1
X_7574_ _1936_ _3070_ _1961_ _3075_ _3237_ VGND 
+ VGND
+ VPWR VPWR _3238_ sky130_fd_sc_hd__o221a_1
X_7575_ _2015_ _3089_ _1972_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3239_ sky130_fd_sc_hd__o22a_1
X_7576_ _1965_ _3085_ _1998_ _3087_ _3239_ VGND 
+ VGND
+ VPWR VPWR _3240_ sky130_fd_sc_hd__o221a_1
X_7577_ _1983_ _3097_ _1959_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3241_ sky130_fd_sc_hd__o22a_1
X_7578_ _1954_ _3104_ _1952_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3242_ sky130_fd_sc_hd__o22a_1
X_7579_ _2007_ _3100_ _1982_ _3102_ _3242_ VGND 
+ VGND
+ VPWR VPWR _3243_ sky130_fd_sc_hd__o221a_1
X_7580_ _2001_ _3095_ _3241_ _3243_ VGND VGND 
+ VPWR
+ VPWR _3244_ sky130_fd_sc_hd__o211a_1
X_7581_ _2008_ _3115_ _1948_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3245_ sky130_fd_sc_hd__o22a_1
X_7582_ _1966_ _3111_ _1978_ _3113_ _3245_ VGND 
+ VGND
+ VPWR VPWR _3246_ sky130_fd_sc_hd__o221a_1
X_7583_ _1938_ _3125_ _1941_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3247_ sky130_fd_sc_hd__o22a_1
X_7584_ _1958_ _3121_ _1943_ _3123_ _3247_ VGND 
+ VGND
+ VPWR VPWR _3248_ sky130_fd_sc_hd__o221a_1
X_7585_ _1967_ _3135_ _1944_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3249_ sky130_fd_sc_hd__o22a_1
X_7586_ _1977_ _3131_ _1951_ _3133_ _3249_ VGND 
+ VGND
+ VPWR VPWR _3250_ sky130_fd_sc_hd__o221a_1
X_7587_ _1971_ _3145_ _1962_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3251_ sky130_fd_sc_hd__o22a_1
X_7588_ _1995_ _3141_ _1964_ _3143_ _3251_ VGND 
+ VGND
+ VPWR VPWR _3252_ sky130_fd_sc_hd__o221a_1
X_7589_ _3246_ _3248_ _3250_ _3252_ VGND VGND 
+ VPWR
+ VPWR _3253_ sky130_fd_sc_hd__and4_1
X_7590_ _3238_ _3240_ _3244_ _3253_ VGND VGND 
+ VPWR
+ VPWR _0140_ sky130_fd_sc_hd__nand4_4
X_7591_ _1866_ _3078_ _1847_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3254_ sky130_fd_sc_hd__o22a_1
X_7592_ _1879_ _3070_ _1925_ _3075_ _3254_ VGND 
+ VGND
+ VPWR VPWR _3255_ sky130_fd_sc_hd__o221a_1
X_7593_ _1917_ _3089_ _1904_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3256_ sky130_fd_sc_hd__o22a_1
X_7594_ _1914_ _3085_ _1908_ _3087_ _3256_ VGND 
+ VGND
+ VPWR VPWR _3257_ sky130_fd_sc_hd__o221a_1
X_7595_ _1860_ _3097_ _1927_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3258_ sky130_fd_sc_hd__o22a_1
X_7596_ _1897_ _3104_ _1898_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3259_ sky130_fd_sc_hd__o22a_1
X_7597_ _1911_ _3100_ _1871_ _3102_ _3259_ VGND 
+ VGND
+ VPWR VPWR _3260_ sky130_fd_sc_hd__o221a_1
X_7598_ _1915_ _3095_ _3258_ _3260_ VGND VGND 
+ VPWR
+ VPWR _3261_ sky130_fd_sc_hd__o211a_1
X_7599_ _1862_ _3115_ _1878_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3262_ sky130_fd_sc_hd__o22a_1
X_7600_ _1910_ _3111_ _1902_ _3113_ _3262_ VGND 
+ VGND
+ VPWR VPWR _3263_ sky130_fd_sc_hd__o221a_1
X_7601_ _1886_ _3125_ _1850_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3264_ sky130_fd_sc_hd__o22a_1
X_7602_ _1926_ _3121_ _1901_ _3123_ _3264_ VGND 
+ VGND
+ VPWR VPWR _3265_ sky130_fd_sc_hd__o221a_1
X_7603_ _1909_ _3135_ _1861_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3266_ sky130_fd_sc_hd__o22a_1
X_7604_ _1853_ _3131_ _1867_ _3133_ _3266_ VGND 
+ VGND
+ VPWR VPWR _3267_ sky130_fd_sc_hd__o221a_1
X_7605_ _1892_ _3145_ _1854_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3268_ sky130_fd_sc_hd__o22a_1
X_7606_ _1916_ _3141_ _1924_ _3143_ _3268_ VGND 
+ VGND
+ VPWR VPWR _3269_ sky130_fd_sc_hd__o221a_1
X_7607_ _3263_ _3265_ _3267_ _3269_ VGND VGND 
+ VPWR
+ VPWR _3270_ sky130_fd_sc_hd__and4_1
X_7608_ _3255_ _3257_ _3261_ _3270_ VGND VGND 
+ VPWR
+ VPWR _0142_ sky130_fd_sc_hd__nand4_4
X_7609_ _1401_ _3078_ _1169_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3271_ sky130_fd_sc_hd__o22a_1
X_7610_ _1397_ _3070_ _1207_ _3075_ _3271_ VGND 
+ VGND
+ VPWR VPWR _3272_ sky130_fd_sc_hd__o221a_1
X_7611_ _1156_ _3089_ _1287_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3273_ sky130_fd_sc_hd__o22a_1
X_7612_ _1191_ _3085_ _1263_ _3087_ _3273_ VGND 
+ VGND
+ VPWR VPWR _3274_ sky130_fd_sc_hd__o221a_1
X_7613_ _1336_ _3097_ _1197_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3275_ sky130_fd_sc_hd__o22a_2
X_7614_ _1279_ _3104_ _1407_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3276_ sky130_fd_sc_hd__o22a_1
X_7615_ _1254_ _3100_ _1314_ _3102_ _3276_ VGND 
+ VGND
+ VPWR VPWR _3277_ sky130_fd_sc_hd__o221a_1
X_7616_ _1244_ _3095_ _3275_ _3277_ VGND VGND 
+ VPWR
+ VPWR _3278_ sky130_fd_sc_hd__o211a_1
X_7617_ _1326_ _3115_ _1395_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3279_ sky130_fd_sc_hd__o22a_1
X_7618_ _1201_ _3111_ _1343_ _3113_ _3279_ VGND 
+ VGND
+ VPWR VPWR _3280_ sky130_fd_sc_hd__o221a_1
X_7619_ _1139_ _3125_ _1301_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3281_ sky130_fd_sc_hd__o22a_1
X_7620_ _1240_ _3121_ _1376_ _3123_ _3281_ VGND 
+ VGND
+ VPWR VPWR _3282_ sky130_fd_sc_hd__o221a_1
X_7621_ _1164_ _3135_ _1365_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3283_ sky130_fd_sc_hd__o22a_1
X_7622_ _1173_ _3131_ _1360_ _3133_ _3283_ VGND 
+ VGND
+ VPWR VPWR _3284_ sky130_fd_sc_hd__o221a_1
X_7623_ _1359_ _3145_ _1185_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3285_ sky130_fd_sc_hd__o22a_1
X_7624_ _1178_ _3141_ _1189_ _3143_ _3285_ VGND 
+ VGND
+ VPWR VPWR _3286_ sky130_fd_sc_hd__o221a_1
X_7625_ _3280_ _3282_ _3284_ _3286_ VGND VGND 
+ VPWR
+ VPWR _3287_ sky130_fd_sc_hd__and4_1
X_7626_ _3272_ _3274_ _3278_ _3287_ VGND VGND 
+ VPWR
+ VPWR _0144_ sky130_fd_sc_hd__nand4_4
X_7627_ _2601_ _3078_ _2637_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3288_ sky130_fd_sc_hd__o22a_1
X_7628_ _2536_ _3070_ _2662_ _3075_ _3288_ VGND 
+ VGND
+ VPWR VPWR _3289_ sky130_fd_sc_hd__o221a_1
X_7629_ _2675_ _3089_ _2603_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3290_ sky130_fd_sc_hd__o22a_1
X_7630_ _2667_ _3085_ _2535_ _3087_ _3290_ VGND 
+ VGND
+ VPWR VPWR _3291_ sky130_fd_sc_hd__o221a_1
X_7631_ _2591_ _3097_ _2673_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3292_ sky130_fd_sc_hd__o22a_1
X_7632_ _2609_ _3104_ _2578_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3293_ sky130_fd_sc_hd__o22a_1
X_7633_ _2657_ _3100_ _2540_ _3102_ _3293_ VGND 
+ VGND
+ VPWR VPWR _3294_ sky130_fd_sc_hd__o221a_1
X_7634_ _2664_ _3095_ _3292_ _3294_ VGND VGND 
+ VPWR
+ VPWR _3295_ sky130_fd_sc_hd__o211a_1
X_7635_ _2602_ _3115_ _2607_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3296_ sky130_fd_sc_hd__o22a_1
X_7636_ _2670_ _3111_ _2559_ _3113_ _3296_ VGND 
+ VGND
+ VPWR VPWR _3297_ sky130_fd_sc_hd__o221a_1
X_7637_ _2633_ _3125_ _2568_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3298_ sky130_fd_sc_hd__o22a_1
X_7638_ _2618_ _3121_ _2608_ _3123_ _3298_ VGND 
+ VGND
+ VPWR VPWR _3299_ sky130_fd_sc_hd__o221a_1
X_7639_ _2632_ _3135_ _2583_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3300_ sky130_fd_sc_hd__o22a_1
X_7640_ _2644_ _3131_ _2580_ _3133_ _3300_ VGND 
+ VGND
+ VPWR VPWR _3301_ sky130_fd_sc_hd__o221a_1
X_7641_ _2547_ _3145_ _2663_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3302_ sky130_fd_sc_hd__o22a_1
X_7642_ _2631_ _3141_ _2669_ _3143_ _3302_ VGND 
+ VGND
+ VPWR VPWR _3303_ sky130_fd_sc_hd__o221a_1
X_7643_ _3297_ _3299_ _3301_ _3303_ VGND VGND 
+ VPWR
+ VPWR _3304_ sky130_fd_sc_hd__and4_1
X_7644_ _3289_ _3291_ _3295_ _3304_ VGND VGND 
+ VPWR
+ VPWR _0146_ sky130_fd_sc_hd__nand4_4
X_7645_ _2466_ _3078_ _2422_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3305_ sky130_fd_sc_hd__o22a_1
X_7646_ _2455_ _3070_ _2382_ _3075_ _3305_ VGND 
+ VGND
+ VPWR VPWR _3306_ sky130_fd_sc_hd__o221a_2
X_7647_ _2469_ _3089_ _2499_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3307_ sky130_fd_sc_hd__o22a_1
X_7648_ _2377_ _3085_ _2509_ _3087_ _3307_ VGND 
+ VGND
+ VPWR VPWR _3308_ sky130_fd_sc_hd__o221a_1
X_7649_ _2449_ _3097_ _2369_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3309_ sky130_fd_sc_hd__o22a_2
X_7650_ _2516_ _3104_ _2517_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3310_ sky130_fd_sc_hd__o22a_1
X_7651_ _2480_ _3100_ _2462_ _3102_ _3310_ VGND 
+ VGND
+ VPWR VPWR _3311_ sky130_fd_sc_hd__o221a_1
X_7652_ _2468_ _3095_ _3309_ _3311_ VGND VGND 
+ VPWR
+ VPWR _3312_ sky130_fd_sc_hd__o211a_1
X_7653_ _2432_ _3115_ _2437_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3313_ sky130_fd_sc_hd__o22a_1
X_7654_ _2375_ _3111_ _2442_ _3113_ _3313_ VGND 
+ VGND
+ VPWR VPWR _3314_ sky130_fd_sc_hd__o221a_1
X_7655_ _2399_ _3125_ _2482_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3315_ sky130_fd_sc_hd__o22a_1
X_7656_ _2419_ _3121_ _2460_ _3123_ _3315_ VGND 
+ VGND
+ VPWR VPWR _3316_ sky130_fd_sc_hd__o221a_1
X_7657_ _2383_ _3135_ _2467_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3317_ sky130_fd_sc_hd__o22a_1
X_7658_ _2411_ _3131_ _2448_ _3133_ _3317_ VGND 
+ VGND
+ VPWR VPWR _3318_ sky130_fd_sc_hd__o221a_1
X_7659_ _2389_ _3145_ _2371_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3319_ sky130_fd_sc_hd__o22a_1
X_7660_ _2487_ _3141_ _2400_ _3143_ _3319_ VGND 
+ VGND
+ VPWR VPWR _3320_ sky130_fd_sc_hd__o221a_1
X_7661_ _3314_ _3316_ _3318_ _3320_ VGND VGND 
+ VPWR
+ VPWR _3321_ sky130_fd_sc_hd__and4_2
X_7662_ _3306_ _3308_ _3312_ _3321_ VGND VGND 
+ VPWR
+ VPWR _0148_ sky130_fd_sc_hd__nand4_4
X_7663_ _2337_ _3078_ _2289_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3322_ sky130_fd_sc_hd__o22a_1
X_7664_ _2312_ _3070_ _2265_ _3075_ _3322_ VGND 
+ VGND
+ VPWR VPWR _3323_ sky130_fd_sc_hd__o221a_2
X_7665_ _2292_ _3089_ _2353_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3324_ sky130_fd_sc_hd__o22a_1
X_7666_ _2331_ _3085_ _2297_ _3087_ _3324_ VGND 
+ VGND
+ VPWR VPWR _3325_ sky130_fd_sc_hd__o221a_1
X_7667_ _2301_ _3097_ _2258_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3326_ sky130_fd_sc_hd__o22a_1
X_7668_ _2350_ _3104_ _2349_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3327_ sky130_fd_sc_hd__o22a_1
X_7669_ _2254_ _3100_ _2344_ _3102_ _3327_ VGND 
+ VGND
+ VPWR VPWR _3328_ sky130_fd_sc_hd__o221a_1
X_7670_ _2279_ _3095_ _3326_ _3328_ VGND VGND 
+ VPWR
+ VPWR _3329_ sky130_fd_sc_hd__o211a_1
X_7671_ _2354_ _3115_ _2336_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3330_ sky130_fd_sc_hd__o22a_1
X_7672_ _2253_ _3111_ _2357_ _3113_ _3330_ VGND 
+ VGND
+ VPWR VPWR _3331_ sky130_fd_sc_hd__o221a_1
X_7673_ _2275_ _3125_ _2308_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3332_ sky130_fd_sc_hd__o22a_1
X_7674_ _2271_ _3121_ _2313_ _3123_ _3332_ VGND 
+ VGND
+ VPWR VPWR _3333_ sky130_fd_sc_hd__o221a_1
X_7675_ _2266_ _3135_ _2327_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3334_ sky130_fd_sc_hd__o22a_1
X_7676_ _2259_ _3131_ _2307_ _3133_ _3334_ VGND 
+ VGND
+ VPWR VPWR _3335_ sky130_fd_sc_hd__o221a_1
X_7677_ _2306_ _3145_ _2276_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3336_ sky130_fd_sc_hd__o22a_1
X_7678_ _2288_ _3141_ _2264_ _3143_ _3336_ VGND 
+ VGND
+ VPWR VPWR _3337_ sky130_fd_sc_hd__o221a_1
X_7679_ _3331_ _3333_ _3335_ _3337_ VGND VGND 
+ VPWR
+ VPWR _3338_ sky130_fd_sc_hd__and4_2
X_7680_ _3323_ _3325_ _3329_ _3338_ VGND VGND 
+ VPWR
+ VPWR _0150_ sky130_fd_sc_hd__nand4_4
X_7681_ _2177_ _3078_ _2196_ _3080_ VGND VGND 
+ VPWR
+ VPWR _3339_ sky130_fd_sc_hd__o22a_1
X_7682_ _2202_ _3070_ _2140_ _3075_ _3339_ VGND 
+ VGND
+ VPWR VPWR _3340_ sky130_fd_sc_hd__o221a_1
X_7683_ _2242_ _3089_ _2119_ _3091_ VGND VGND 
+ VPWR
+ VPWR _3341_ sky130_fd_sc_hd__o22a_1
X_7684_ _2151_ _3085_ _2194_ _3087_ _3341_ VGND 
+ VGND
+ VPWR VPWR _3342_ sky130_fd_sc_hd__o221a_1
X_7685_ _2169_ _3097_ _2139_ _1697_ VGND VGND 
+ VPWR
+ VPWR _3343_ sky130_fd_sc_hd__o22a_1
X_7686_ _2108_ _3104_ _2125_ _3106_ VGND VGND 
+ VPWR
+ VPWR _3344_ sky130_fd_sc_hd__o22a_1
X_7687_ _2109_ _3100_ _2190_ _3102_ _3344_ VGND 
+ VGND
+ VPWR VPWR _3345_ sky130_fd_sc_hd__o221a_1
X_7688_ _2236_ _3095_ _3343_ _3345_ VGND VGND 
+ VPWR
+ VPWR _3346_ sky130_fd_sc_hd__o211a_1
X_7689_ _2187_ _3115_ _2182_ _3117_ VGND VGND 
+ VPWR
+ VPWR _3347_ sky130_fd_sc_hd__o22a_1
X_7690_ _2152_ _3111_ _2165_ _3113_ _3347_ VGND 
+ VGND
+ VPWR VPWR _3348_ sky130_fd_sc_hd__o221a_1
X_7691_ _2141_ _3125_ _2223_ _3127_ VGND VGND 
+ VPWR
+ VPWR _3349_ sky130_fd_sc_hd__o22a_1
X_7692_ _2245_ _3121_ _2126_ _3123_ _3349_ VGND 
+ VGND
+ VPWR VPWR _3350_ sky130_fd_sc_hd__o221a_1
X_7693_ _2147_ _3135_ _2175_ _3137_ VGND VGND 
+ VPWR
+ VPWR _3351_ sky130_fd_sc_hd__o22a_1
X_7694_ _2212_ _3131_ _2118_ _3133_ _3351_ VGND 
+ VGND
+ VPWR VPWR _3352_ sky130_fd_sc_hd__o221a_1
X_7695_ _2207_ _3145_ _2157_ _3147_ VGND VGND 
+ VPWR
+ VPWR _3353_ sky130_fd_sc_hd__o22a_1
X_7696_ _2219_ _3141_ _2156_ _3143_ _3353_ VGND 
+ VGND
+ VPWR VPWR _3354_ sky130_fd_sc_hd__o221a_1
X_7697_ _3348_ _3350_ _3352_ _3354_ VGND VGND 
+ VPWR
+ VPWR _3355_ sky130_fd_sc_hd__and4_1
X_7698_ _3340_ _3342_ _3346_ _3355_ VGND VGND 
+ VPWR
+ VPWR _0152_ sky130_fd_sc_hd__nand4_4
X_7699_ _4413_ VGND VGND VPWR VPWR _3356_ sky130_fd_sc_hd__clkbuf_1
X_7700_ _3356_ VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__clkbuf_1
X_7701_ _4412_ VGND VGND VPWR VPWR _3357_ sky130_fd_sc_hd__clkbuf_1
X_7702_ _3357_ VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__clkbuf_1
X_7703_ _4410_ VGND VGND VPWR VPWR _3358_ sky130_fd_sc_hd__clkbuf_1
X_7704_ _3358_ VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__clkbuf_1
X_7705_ _4409_ VGND VGND VPWR VPWR _3359_ sky130_fd_sc_hd__clkbuf_1
X_7706_ _3359_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__clkbuf_1
X_7707_ \hkspi.state[1]\ \hkspi.state[4]\ VGND VGND VPWR VPWR 
+ _0155_
+ sky130_fd_sc_hd__nor2_1
X_7708_ \hkspi.addr[0]\ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkinv_2
X_7709_ \hkspi.addr[1]\ \hkspi.addr[0]\ VGND VGND VPWR VPWR 
+ _3360_
+ sky130_fd_sc_hd__nand2_1
X_7710_ \hkspi.addr[1]\ \hkspi.addr[0]\ _3360_ VGND VGND VPWR 
+ VPWR
+ _0157_ sky130_fd_sc_hd__o21a_1
X_7711_ _3360_ VGND VGND VPWR VPWR _3361_ sky130_fd_sc_hd__inv_2
X_7712_ \hkspi.addr[2]\ _3361_ \hkspi.addr[2]\ _3361_ VGND VGND 
+ VPWR
+ VPWR _0158_ sky130_fd_sc_hd__o2bb2a_1
X_7713_ \hkspi.addr[2]\ _3361_ \hkspi.addr[3]\ VGND VGND VPWR 
+ VPWR
+ _3362_ sky130_fd_sc_hd__and3_1
X_7714_ \hkspi.addr[2]\ _3361_ \hkspi.addr[3]\ VGND VGND VPWR 
+ VPWR
+ _3363_ sky130_fd_sc_hd__a21oi_1
X_7715_ _3362_ _3363_ VGND VGND VPWR VPWR 
+ _0159_
+ sky130_fd_sc_hd__nor2_1
X_7716_ \hkspi.addr[4]\ _3362_ VGND VGND VPWR VPWR 
+ _3364_
+ sky130_fd_sc_hd__nand2_1
X_7717_ \hkspi.addr[4]\ _3362_ _3364_ VGND VGND VPWR 
+ VPWR
+ _0160_ sky130_fd_sc_hd__o21a_1
X_7718_ _3364_ VGND VGND VPWR VPWR _3365_ sky130_fd_sc_hd__inv_2
X_7719_ \hkspi.addr[5]\ _3365_ VGND VGND VPWR VPWR 
+ _3366_
+ sky130_fd_sc_hd__nand2_1
X_7720_ \hkspi.addr[5]\ _3365_ _3366_ VGND VGND VPWR 
+ VPWR
+ _0161_ sky130_fd_sc_hd__o21a_1
X_7721_ _3366_ VGND VGND VPWR VPWR _3367_ sky130_fd_sc_hd__inv_2
X_7722_ \hkspi.addr[6]\ _3367_ VGND VGND VPWR VPWR 
+ _3368_
+ sky130_fd_sc_hd__nand2_1
X_7723_ \hkspi.addr[6]\ _3367_ _3368_ VGND VGND VPWR 
+ VPWR
+ _0162_ sky130_fd_sc_hd__o21a_1
X_7724_ \hkspi.addr[7]\ VGND VGND VPWR VPWR _3369_ sky130_fd_sc_hd__inv_2
X_7725_ \hkspi.addr[6]\ _3367_ _3369_ \hkspi.addr[7]\ _3368_ VGND 
+ VGND
+ VPWR VPWR _0163_ sky130_fd_sc_hd__a32o_1
X_7726_ \hkspi.fixed[0]\ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkinv_4
X_7727_ \hkspi.fixed[1]\ VGND VGND VPWR VPWR _3370_ sky130_fd_sc_hd__inv_2
X_7728_ _3370_ _0164_ \hkspi.fixed[1]\ \hkspi.fixed[0]\ VGND VGND 
+ VPWR
+ VPWR _0165_ sky130_fd_sc_hd__a22o_1
X_7729_ _3370_ _0164_ \hkspi.fixed[2]\ VGND VGND VPWR 
+ VPWR
+ _3371_ sky130_fd_sc_hd__a21oi_1
X_7730_ _3370_ _0164_ \hkspi.fixed[2]\ _3371_ VGND VGND 
+ VPWR
+ VPWR _0166_ sky130_fd_sc_hd__a31oi_1
X_7731_ _1080_ _0169_ VGND VGND VPWR VPWR 
+ _3372_
+ sky130_fd_sc_hd__and2_1
X_7732_ _3372_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_7733_ net199 net202 \wbbd_state[7]\ VGND VGND VPWR 
+ VPWR
+ _3373_ sky130_fd_sc_hd__and3_1
X_7734_ net202 net200 \wbbd_state[9]\ VGND VGND VPWR 
+ VPWR
+ _3374_ sky130_fd_sc_hd__and3_1
X_7735_ \wbbd_state[8]\ _1472_ _3373_ _3374_ VGND VGND 
+ VPWR
+ VPWR _0168_ sky130_fd_sc_hd__a211o_1
X_7736_ \wbbd_state[7]\ net171 VGND VGND VPWR VPWR 
+ _3375_
+ sky130_fd_sc_hd__and2_1
X_7737_ \wbbd_state[9]\ net180 \wbbd_state[8]\ net194 _3375_ VGND 
+ VGND
+ VPWR VPWR _0170_ sky130_fd_sc_hd__a221o_1
X_7738_ \wbbd_state[7]\ net172 VGND VGND VPWR VPWR 
+ _3376_
+ sky130_fd_sc_hd__and2_1
X_7739_ \wbbd_state[9]\ net181 \wbbd_state[8]\ net195 _3376_ VGND 
+ VGND
+ VPWR VPWR _0171_ sky130_fd_sc_hd__a221o_1
X_7740_ \wbbd_state[7]\ net173 VGND VGND VPWR VPWR 
+ _3377_
+ sky130_fd_sc_hd__and2_1
X_7741_ \wbbd_state[9]\ net182 \wbbd_state[8]\ net165 _3377_ VGND 
+ VGND
+ VPWR VPWR _0172_ sky130_fd_sc_hd__a221o_1
X_7742_ \wbbd_state[7]\ net174 VGND VGND VPWR VPWR 
+ _3378_
+ sky130_fd_sc_hd__and2_1
X_7743_ \wbbd_state[9]\ net183 \wbbd_state[8]\ net166 _3378_ VGND 
+ VGND
+ VPWR VPWR _0173_ sky130_fd_sc_hd__a221o_1
X_7744_ \wbbd_state[7]\ net176 VGND VGND VPWR VPWR 
+ _3379_
+ sky130_fd_sc_hd__and2_1
X_7745_ \wbbd_state[9]\ net184 \wbbd_state[8]\ net167 _3379_ VGND 
+ VGND
+ VPWR VPWR _0174_ sky130_fd_sc_hd__a221o_1
X_7746_ \wbbd_state[7]\ net177 VGND VGND VPWR VPWR 
+ _3380_
+ sky130_fd_sc_hd__and2_1
X_7747_ \wbbd_state[9]\ net185 \wbbd_state[8]\ net168 _3380_ VGND 
+ VGND
+ VPWR VPWR _0175_ sky130_fd_sc_hd__a221o_1
X_7748_ \wbbd_state[7]\ net178 VGND VGND VPWR VPWR 
+ _3381_
+ sky130_fd_sc_hd__and2_1
X_7749_ \wbbd_state[9]\ net187 \wbbd_state[8]\ net169 _3381_ VGND 
+ VGND
+ VPWR VPWR _0176_ sky130_fd_sc_hd__a221o_1
X_7750_ \wbbd_state[7]\ net179 VGND VGND VPWR VPWR 
+ _3382_
+ sky130_fd_sc_hd__and2_1
X_7751_ \wbbd_state[9]\ net188 \wbbd_state[8]\ net170 _3382_ VGND 
+ VGND
+ VPWR VPWR _0177_ sky130_fd_sc_hd__a221o_1
X_7752_ net153 VGND VGND VPWR VPWR _3383_ sky130_fd_sc_hd__inv_2
X_7753_ net142 net131 VGND VGND VPWR VPWR 
+ _3384_
+ sky130_fd_sc_hd__or2_2
X_7754_ net156 _3383_ _3384_ VGND VGND VPWR 
+ VPWR
+ _3385_ sky130_fd_sc_hd__or3_4
X_7755_ _3385_ VGND VGND VPWR VPWR _3386_ sky130_fd_sc_hd__inv_2
X_7756_ net144 _1795_ _1791_ VGND VGND VPWR 
+ VPWR
+ _3387_ sky130_fd_sc_hd__or3_1
X_7757_ _3387_ VGND VGND VPWR VPWR _3388_ sky130_fd_sc_hd__buf_4
X_7758_ _3388_ VGND VGND VPWR VPWR _3389_ sky130_fd_sc_hd__clkinv_2
X_7759_ net158 net157 net159 net160 VGND VGND 
+ VPWR
+ VPWR _3390_ sky130_fd_sc_hd__or4_4
X_7760_ _3390_ VGND VGND VPWR VPWR _3391_ sky130_fd_sc_hd__inv_2
X_7761_ _3386_ _3389_ _3391_ VGND VGND VPWR 
+ VPWR
+ _3392_ sky130_fd_sc_hd__and3_2
X_7762_ net156 VGND VGND VPWR VPWR _3393_ sky130_fd_sc_hd__clkinv_4
X_7763_ _3393_ net153 _3384_ VGND VGND VPWR 
+ VPWR
+ _3394_ sky130_fd_sc_hd__or3_1
X_7764_ _3394_ VGND VGND VPWR VPWR _3395_ sky130_fd_sc_hd__clkbuf_16
X_7765_ net157 VGND VGND VPWR VPWR _3396_ sky130_fd_sc_hd__inv_6
X_7766_ _3384_ VGND VGND VPWR VPWR _3397_ sky130_fd_sc_hd__inv_2
X_7767_ _3393_ _3383_ _3397_ VGND VGND VPWR 
+ VPWR
+ _3398_ sky130_fd_sc_hd__or3_2
X_7768_ net139 net138 net141 net140 VGND VGND 
+ VPWR
+ VPWR _3399_ sky130_fd_sc_hd__nand4_1
X_7769_ net160 VGND VGND VPWR VPWR _3400_ sky130_fd_sc_hd__clkinv_4
X_7770_ net137 net136 VGND VGND VPWR VPWR 
+ _3401_
+ sky130_fd_sc_hd__nand2_1
X_7771_ net133 net132 net135 net134 VGND VGND 
+ VPWR
+ VPWR _3402_ sky130_fd_sc_hd__nand4_1
X_7772_ net159 VGND VGND VPWR VPWR _3403_ sky130_fd_sc_hd__inv_2
X_7773_ net158 VGND VGND VPWR VPWR _3404_ sky130_fd_sc_hd__inv_6
X_7774_ _3403_ _3404_ net162 net161 VGND VGND 
+ VPWR
+ VPWR _3405_ sky130_fd_sc_hd__nand4bb_1
X_7775_ _3400_ _3401_ _3402_ _3405_ VGND VGND 
+ VPWR
+ VPWR _3406_ sky130_fd_sc_hd__or4_1
X_7776_ _3396_ _3398_ _3399_ _3406_ VGND VGND 
+ VPWR
+ VPWR _3407_ sky130_fd_sc_hd__or4_1
X_7777_ _3407_ VGND VGND VPWR VPWR _3408_ sky130_fd_sc_hd__inv_2
X_7778_ _1795_ _3408_ net143 _3407_ VGND VGND 
+ VPWR
+ VPWR _3409_ sky130_fd_sc_hd__o22a_1
X_7779_ net144 net143 _1796_ VGND VGND VPWR 
+ VPWR
+ _3410_ sky130_fd_sc_hd__o21ai_2
X_7780_ _3410_ VGND VGND VPWR VPWR _3411_ sky130_fd_sc_hd__inv_2
X_7781_ net146 net145 VGND VGND VPWR VPWR 
+ _3412_
+ sky130_fd_sc_hd__nand2_1
X_7782_ net144 net143 _3412_ _1791_ _1796_ VGND 
+ VGND
+ VPWR VPWR _3413_ sky130_fd_sc_hd__a32o_2
X_7783_ _3411_ _3408_ net144 _3407_ _3413_ VGND 
+ VGND
+ VPWR VPWR _3414_ sky130_fd_sc_hd__a221o_1
X_7784_ _3409_ _3414_ VGND VGND VPWR VPWR 
+ _3415_
+ sky130_fd_sc_hd__or2_1
X_7785_ _3404_ _3396_ _3398_ VGND VGND VPWR 
+ VPWR
+ _3416_ sky130_fd_sc_hd__or3_1
X_7786_ _3416_ VGND VGND VPWR VPWR _3417_ sky130_fd_sc_hd__inv_2
X_7787_ _3403_ _3416_ VGND VGND VPWR VPWR 
+ _3418_
+ sky130_fd_sc_hd__or2_1
X_7788_ net159 _3417_ _3418_ VGND VGND VPWR 
+ VPWR
+ _3419_ sky130_fd_sc_hd__o21ai_2
X_7789_ net159 _3417_ net160 _3400_ _3418_ VGND 
+ VGND
+ VPWR VPWR _3420_ sky130_fd_sc_hd__a32o_1
X_7790_ _3419_ _3420_ VGND VGND VPWR VPWR 
+ _3421_
+ sky130_fd_sc_hd__nand2_1
X_7791_ _3396_ _3398_ VGND VGND VPWR VPWR 
+ _3422_
+ sky130_fd_sc_hd__nor2_1
X_7792_ net158 _3422_ VGND VGND VPWR VPWR 
+ _3423_
+ sky130_fd_sc_hd__nor2_1
X_7793_ _3396_ _3398_ _3422_ VGND VGND VPWR 
+ VPWR
+ _3424_ sky130_fd_sc_hd__a21o_2
X_7794_ _3417_ _3423_ _3424_ VGND VGND VPWR 
+ VPWR
+ _3425_ sky130_fd_sc_hd__o21ai_2
X_7795_ _3421_ _3425_ VGND VGND VPWR VPWR 
+ _3426_
+ sky130_fd_sc_hd__or2_2
X_7796_ _3415_ _3426_ VGND VGND VPWR VPWR 
+ _3427_
+ sky130_fd_sc_hd__or2_1
X_7797_ _3427_ VGND VGND VPWR VPWR _3428_ sky130_fd_sc_hd__buf_2
X_7798_ _3395_ _3428_ VGND VGND VPWR VPWR 
+ _3429_
+ sky130_fd_sc_hd__nor2_2
X_7799_ net142 VGND VGND VPWR VPWR _3430_ sky130_fd_sc_hd__inv_6
X_7800_ _3430_ net131 net156 VGND VGND VPWR 
+ VPWR
+ _3431_ sky130_fd_sc_hd__or3_4
X_7801_ _3383_ _3431_ VGND VGND VPWR VPWR 
+ _3432_
+ sky130_fd_sc_hd__or2_1
X_7802_ _3432_ VGND VGND VPWR VPWR _3433_ sky130_fd_sc_hd__buf_6
X_7803_ _3428_ _3433_ VGND VGND VPWR VPWR 
+ _3434_
+ sky130_fd_sc_hd__nor2_1
X_7804_ _3430_ _3393_ net153 VGND VGND VPWR 
+ VPWR
+ _3435_ sky130_fd_sc_hd__or3_4
X_7805_ net131 _3435_ VGND VGND VPWR VPWR 
+ _3436_
+ sky130_fd_sc_hd__or2_1
X_7806_ _3436_ VGND VGND VPWR VPWR _3437_ sky130_fd_sc_hd__buf_8
X_7807_ _3390_ _3437_ VGND VGND VPWR VPWR 
+ _3438_
+ sky130_fd_sc_hd__or2_2
X_7808_ _3388_ _3438_ VGND VGND VPWR VPWR 
+ _3439_
+ sky130_fd_sc_hd__nor2_2
X_7809_ net159 net160 net158 _3396_ VGND VGND 
+ VPWR
+ VPWR _3440_ sky130_fd_sc_hd__or4_1
X_7810_ _3388_ _3440_ VGND VGND VPWR VPWR 
+ _3441_
+ sky130_fd_sc_hd__or2_1
X_7811_ _3441_ VGND VGND VPWR VPWR _3442_ sky130_fd_sc_hd__clkbuf_8
X_7812_ net156 net153 _3384_ VGND VGND VPWR 
+ VPWR
+ _3443_ sky130_fd_sc_hd__or3_1
X_7813_ _3443_ VGND VGND VPWR VPWR _3444_ sky130_fd_sc_hd__clkbuf_16
X_7814_ _3430_ net131 _3393_ _3383_ VGND VGND 
+ VPWR
+ VPWR _3445_ sky130_fd_sc_hd__or4_1
X_7815_ _3445_ VGND VGND VPWR VPWR _3446_ sky130_fd_sc_hd__buf_12
X_7816_ _3442_ _3446_ VGND VGND VPWR VPWR 
+ _3447_
+ sky130_fd_sc_hd__or2_1
X_7817_ _3444_ VGND VGND VPWR VPWR _3448_ sky130_fd_sc_hd__inv_2
X_7818_ net159 net160 _3404_ net157 VGND VGND 
+ VPWR
+ VPWR _3449_ sky130_fd_sc_hd__or4_1
X_7819_ _3449_ VGND VGND VPWR VPWR _3450_ sky130_fd_sc_hd__clkbuf_4
X_7820_ _3450_ VGND VGND VPWR VPWR _3451_ sky130_fd_sc_hd__inv_2
X_7821_ _3393_ _3383_ _3384_ VGND VGND VPWR 
+ VPWR
+ _3452_ sky130_fd_sc_hd__or3_4
X_7822_ _3442_ _3452_ VGND VGND VPWR VPWR 
+ _3453_
+ sky130_fd_sc_hd__nor2_4
X_7823_ _3417_ _3423_ _3424_ VGND VGND VPWR 
+ VPWR
+ _3454_ sky130_fd_sc_hd__or3b_1
X_7824_ _3421_ _3454_ _3415_ VGND VGND VPWR 
+ VPWR
+ _3455_ sky130_fd_sc_hd__or3_1
X_7825_ _3455_ VGND VGND VPWR VPWR _3456_ sky130_fd_sc_hd__buf_2
X_7826_ _3456_ _3452_ VGND VGND VPWR VPWR 
+ _3457_
+ sky130_fd_sc_hd__or2_1
X_7827_ _3457_ VGND VGND VPWR VPWR _3458_ sky130_fd_sc_hd__inv_2
X_7828_ _3446_ _3450_ _3388_ VGND VGND VPWR 
+ VPWR
+ _3459_ sky130_fd_sc_hd__or3_1
X_7829_ _3459_ VGND VGND VPWR VPWR _3460_ sky130_fd_sc_hd__inv_2
X_7830_ net159 net160 _3404_ _3396_ VGND VGND 
+ VPWR
+ VPWR _3461_ sky130_fd_sc_hd__or4_4
X_7831_ _3461_ VGND VGND VPWR VPWR _3462_ sky130_fd_sc_hd__inv_2
X_7832_ net144 net143 _1791_ VGND VGND VPWR 
+ VPWR
+ _3463_ sky130_fd_sc_hd__or3_1
X_7833_ _3463_ VGND VGND VPWR VPWR _3464_ sky130_fd_sc_hd__buf_8
X_7834_ _3464_ VGND VGND VPWR VPWR _3465_ sky130_fd_sc_hd__clkbuf_16
X_7835_ _3465_ VGND VGND VPWR VPWR _3466_ sky130_fd_sc_hd__inv_4
X_7836_ _3391_ _3466_ _3448_ VGND VGND VPWR 
+ VPWR
+ _3467_ sky130_fd_sc_hd__and3_1
X_7837_ _1794_ net143 _1791_ VGND VGND VPWR 
+ VPWR
+ _3468_ sky130_fd_sc_hd__or3_4
X_7838_ net156 _3384_ _3390_ _3468_ VGND VGND 
+ VPWR
+ VPWR _3469_ sky130_fd_sc_hd__or4_1
X_7839_ net131 VGND VGND VPWR VPWR _3470_ sky130_fd_sc_hd__inv_2
X_7840_ net156 _3383_ net142 _3470_ VGND VGND 
+ VPWR
+ VPWR _3471_ sky130_fd_sc_hd__or4_1
X_7841_ _3471_ VGND VGND VPWR VPWR _3472_ sky130_fd_sc_hd__buf_12
X_7842_ _3450_ _3465_ VGND VGND VPWR VPWR 
+ _3473_
+ sky130_fd_sc_hd__or2_2
X_7843_ _3472_ _3473_ VGND VGND VPWR VPWR 
+ _3474_
+ sky130_fd_sc_hd__or2_2
X_7844_ _3393_ net153 net142 _3470_ VGND VGND 
+ VPWR
+ VPWR _3475_ sky130_fd_sc_hd__or4_1
X_7845_ _3475_ VGND VGND VPWR VPWR _3476_ sky130_fd_sc_hd__buf_8
X_7846_ _3393_ _3383_ net142 _3470_ VGND VGND 
+ VPWR
+ VPWR _3477_ sky130_fd_sc_hd__or4_1
X_7847_ _3477_ VGND VGND VPWR VPWR _3478_ sky130_fd_sc_hd__buf_12
X_7848_ _3473_ _3478_ VGND VGND VPWR VPWR 
+ _3479_
+ sky130_fd_sc_hd__or2_1
X_7849_ net156 net153 net142 _3470_ VGND VGND 
+ VPWR
+ VPWR _3480_ sky130_fd_sc_hd__or4_1
X_7850_ _3480_ VGND VGND VPWR VPWR _3481_ sky130_fd_sc_hd__buf_12
X_7851_ _3461_ _3465_ VGND VGND VPWR VPWR 
+ _3482_
+ sky130_fd_sc_hd__or2_1
X_7852_ _3482_ VGND VGND VPWR VPWR _3483_ sky130_fd_sc_hd__clkbuf_2
X_7853_ _3481_ _3483_ VGND VGND VPWR VPWR 
+ _3484_
+ sky130_fd_sc_hd__or2_1
X_7854_ _3472_ _3483_ VGND VGND VPWR VPWR 
+ _3485_
+ sky130_fd_sc_hd__nor2_1
X_7855_ _3478_ _3483_ VGND VGND VPWR VPWR 
+ _3486_
+ sky130_fd_sc_hd__nor2_1
X_7856_ net158 net157 _3403_ net160 VGND VGND 
+ VPWR
+ VPWR _3487_ sky130_fd_sc_hd__or4_4
X_7857_ _3465_ _3487_ VGND VGND VPWR VPWR 
+ _3488_
+ sky130_fd_sc_hd__or2_1
X_7858_ _3488_ VGND VGND VPWR VPWR _3489_ sky130_fd_sc_hd__dlymetal6s2s_1
X_7859_ _3481_ _3489_ VGND VGND VPWR VPWR 
+ _3490_
+ sky130_fd_sc_hd__nor2_1
X_7860_ _3472_ _3489_ VGND VGND VPWR VPWR 
+ _3491_
+ sky130_fd_sc_hd__nor2_1
X_7861_ _3476_ VGND VGND VPWR VPWR _3492_ sky130_fd_sc_hd__inv_2
X_7862_ _3487_ VGND VGND VPWR VPWR _3493_ sky130_fd_sc_hd__inv_2
X_7863_ _3465_ _3476_ VGND VGND VPWR VPWR 
+ _3494_
+ sky130_fd_sc_hd__or2_1
X_7864_ _3494_ VGND VGND VPWR VPWR _3495_ sky130_fd_sc_hd__buf_6
X_7865_ _3403_ net160 net158 _3396_ VGND VGND 
+ VPWR
+ VPWR _3496_ sky130_fd_sc_hd__or4_4
X_7866_ _3496_ VGND VGND VPWR VPWR _3497_ sky130_fd_sc_hd__buf_2
X_7867_ _3403_ net160 _3404_ net157 VGND VGND 
+ VPWR
+ VPWR _3498_ sky130_fd_sc_hd__or4_4
X_7868_ _3498_ VGND VGND VPWR VPWR _3499_ sky130_fd_sc_hd__clkbuf_4
X_7869_ _3464_ _3499_ VGND VGND VPWR VPWR 
+ _3500_
+ sky130_fd_sc_hd__or2_1
X_7870_ _3500_ VGND VGND VPWR VPWR _3501_ sky130_fd_sc_hd__clkbuf_4
X_7871_ _3472_ _3501_ VGND VGND VPWR VPWR 
+ _3502_
+ sky130_fd_sc_hd__nor2_2
X_7872_ _3404_ _3396_ _3403_ net160 VGND VGND 
+ VPWR
+ VPWR _3503_ sky130_fd_sc_hd__or4_4
X_7873_ _3503_ VGND VGND VPWR VPWR _3504_ sky130_fd_sc_hd__buf_2
X_7874_ _3504_ _3464_ VGND VGND VPWR VPWR 
+ _3505_
+ sky130_fd_sc_hd__or2_2
X_7875_ net158 net157 net159 _3400_ VGND VGND 
+ VPWR
+ VPWR _3506_ sky130_fd_sc_hd__or4_4
X_7876_ _3464_ _3506_ VGND VGND VPWR VPWR 
+ _3507_
+ sky130_fd_sc_hd__or2_2
X_7877_ _3472_ _3507_ VGND VGND VPWR VPWR 
+ _3508_
+ sky130_fd_sc_hd__or2_2
X_7878_ _3440_ _3444_ VGND VGND VPWR VPWR 
+ _3509_
+ sky130_fd_sc_hd__or2_2
X_7879_ _3468_ _3509_ VGND VGND VPWR VPWR 
+ _3510_
+ sky130_fd_sc_hd__nor2_1
X_7880_ _3390_ _3452_ VGND VGND VPWR VPWR 
+ _3511_
+ sky130_fd_sc_hd__or2_2
X_7881_ _3511_ VGND VGND VPWR VPWR _3512_ sky130_fd_sc_hd__inv_2
X_7882_ _3390_ _3446_ VGND VGND VPWR VPWR 
+ _3513_
+ sky130_fd_sc_hd__or2_4
X_7883_ _3513_ VGND VGND VPWR VPWR _3514_ sky130_fd_sc_hd__inv_2
X_7884_ net159 _3400_ _3404_ VGND VGND VPWR 
+ VPWR
+ _3515_ sky130_fd_sc_hd__or3_2
X_7885_ _3472_ _3515_ VGND VGND VPWR VPWR 
+ _3516_
+ sky130_fd_sc_hd__or2_1
X_7886_ _3512_ _3514_ _3509_ _3516_ VGND VGND 
+ VPWR
+ VPWR _3517_ sky130_fd_sc_hd__or4bb_1
X_7887_ _3466_ _3510_ _3517_ VGND VGND VPWR 
+ VPWR
+ _3518_ sky130_fd_sc_hd__o21ai_2
X_7888_ _3465_ _3481_ VGND VGND VPWR VPWR 
+ _3519_
+ sky130_fd_sc_hd__or2_1
X_7889_ net158 _3396_ net159 _3400_ VGND VGND 
+ VPWR
+ VPWR _3520_ sky130_fd_sc_hd__or4_1
X_7890_ _3520_ VGND VGND VPWR VPWR _3521_ sky130_fd_sc_hd__buf_4
X_7891_ _3519_ _3521_ VGND VGND VPWR VPWR 
+ _3522_
+ sky130_fd_sc_hd__or2_1
X_7892_ _3472_ _3476_ _3465_ _3521_ VGND VGND 
+ VPWR
+ VPWR _3523_ sky130_fd_sc_hd__a211o_1
X_7893_ _3478_ _3507_ _3522_ _3523_ VGND VGND 
+ VPWR
+ VPWR _3524_ sky130_fd_sc_hd__o211a_1
X_7894_ _3404_ net157 net159 _3400_ VGND VGND 
+ VPWR
+ VPWR _3525_ sky130_fd_sc_hd__or4_1
X_7895_ _3525_ VGND VGND VPWR VPWR _3526_ sky130_fd_sc_hd__clkbuf_8
X_7896_ _3519_ _3526_ VGND VGND VPWR VPWR 
+ _3527_
+ sky130_fd_sc_hd__or2_1
X_7897_ _3409_ VGND VGND VPWR VPWR _3528_ sky130_fd_sc_hd__inv_2
X_7898_ _3528_ _3414_ VGND VGND VPWR VPWR 
+ _3529_
+ sky130_fd_sc_hd__or2_4
X_7899_ _3454_ _3529_ VGND VGND VPWR VPWR 
+ _3530_
+ sky130_fd_sc_hd__or2_2
X_7900_ _3420_ _3419_ VGND VGND VPWR VPWR 
+ _3531_
+ sky130_fd_sc_hd__or2b_2
X_7901_ _3530_ _3531_ VGND VGND VPWR VPWR 
+ _3532_
+ sky130_fd_sc_hd__or2_1
X_7902_ _3478_ _3532_ VGND VGND VPWR VPWR 
+ _3533_
+ sky130_fd_sc_hd__or2_1
X_7903_ _3404_ _3396_ net159 _3400_ VGND VGND 
+ VPWR
+ VPWR _3534_ sky130_fd_sc_hd__or4_1
X_7904_ _3534_ VGND VGND VPWR VPWR _3535_ sky130_fd_sc_hd__clkbuf_4
X_7905_ _3465_ _3478_ _3526_ _3519_ _3535_ VGND 
+ VGND
+ VPWR VPWR _3536_ sky130_fd_sc_hd__o32a_1
X_7906_ _3495_ _3515_ _3527_ _3533_ _3536_ VGND 
+ VGND
+ VPWR VPWR _3537_ sky130_fd_sc_hd__o2111a_1
X_7907_ _3495_ _3506_ _3518_ _3524_ _3537_ VGND 
+ VGND
+ VPWR VPWR _3538_ sky130_fd_sc_hd__o2111a_2
X_7908_ _3481_ _3507_ VGND VGND VPWR VPWR 
+ _3539_
+ sky130_fd_sc_hd__or2_1
X_7909_ _3478_ _3505_ _3508_ _3538_ _3539_ VGND 
+ VGND
+ VPWR VPWR _3540_ sky130_fd_sc_hd__o2111a_1
X_7910_ _3472_ _3505_ VGND VGND VPWR VPWR 
+ _3541_
+ sky130_fd_sc_hd__or2_1
X_7911_ _3481_ _3505_ VGND VGND VPWR VPWR 
+ _3542_
+ sky130_fd_sc_hd__or2_1
X_7912_ _3504_ _3495_ _3540_ _3541_ _3542_ VGND 
+ VGND
+ VPWR VPWR _3543_ sky130_fd_sc_hd__o2111a_1
X_7913_ _3478_ _3501_ _3495_ _3499_ _3543_ VGND 
+ VGND
+ VPWR VPWR _3544_ sky130_fd_sc_hd__o221ai_1
X_7914_ _3481_ _3501_ VGND VGND VPWR VPWR 
+ _3545_
+ sky130_fd_sc_hd__nor2_1
X_7915_ _3464_ _3497_ VGND VGND VPWR VPWR 
+ _3546_
+ sky130_fd_sc_hd__or2_1
X_7916_ _3478_ _3546_ VGND VGND VPWR VPWR 
+ _3547_
+ sky130_fd_sc_hd__nor2_1
X_7917_ _3502_ _3544_ _3545_ _3547_ VGND VGND 
+ VPWR
+ VPWR _3548_ sky130_fd_sc_hd__nor4_1
X_7918_ _3472_ _3546_ VGND VGND VPWR VPWR 
+ _3549_
+ sky130_fd_sc_hd__or2_1
X_7919_ _3481_ _3546_ VGND VGND VPWR VPWR 
+ _3550_
+ sky130_fd_sc_hd__or2_1
X_7920_ _3495_ _3497_ _3548_ _3549_ _3550_ VGND 
+ VGND
+ VPWR VPWR _3551_ sky130_fd_sc_hd__o2111a_1
X_7921_ _3478_ _3489_ _3551_ VGND VGND VPWR 
+ VPWR
+ _3552_ sky130_fd_sc_hd__o21ai_1
X_7922_ _3466_ _3492_ _3493_ _3552_ VGND VGND 
+ VPWR
+ VPWR _3553_ sky130_fd_sc_hd__a31o_1
X_7923_ _3491_ _3553_ VGND VGND VPWR VPWR 
+ _3554_
+ sky130_fd_sc_hd__or2_1
X_7924_ _3490_ _3554_ VGND VGND VPWR VPWR 
+ _3555_
+ sky130_fd_sc_hd__or2_1
X_7925_ _3486_ _3555_ VGND VGND VPWR VPWR 
+ _3556_
+ sky130_fd_sc_hd__nor2_1
X_7926_ _3476_ _3483_ _3556_ VGND VGND VPWR 
+ VPWR
+ _3557_ sky130_fd_sc_hd__o21ai_1
X_7927_ _3485_ _3557_ VGND VGND VPWR VPWR 
+ _3558_
+ sky130_fd_sc_hd__nor2_1
X_7928_ _3484_ _3558_ VGND VGND VPWR VPWR 
+ _3559_
+ sky130_fd_sc_hd__and2_1
X_7929_ _3479_ _3559_ VGND VGND VPWR VPWR 
+ _3560_
+ sky130_fd_sc_hd__nand2_1
X_7930_ _3473_ _3476_ _3560_ VGND VGND VPWR 
+ VPWR
+ _3561_ sky130_fd_sc_hd__o21ba_1
X_7931_ _3474_ _3561_ VGND VGND VPWR VPWR 
+ _3562_
+ sky130_fd_sc_hd__and2_1
X_7932_ _3383_ _3469_ _3562_ VGND VGND VPWR 
+ VPWR
+ _3563_ sky130_fd_sc_hd__o21ai_1
X_7933_ _3467_ _3563_ VGND VGND VPWR VPWR 
+ _3564_
+ sky130_fd_sc_hd__or2_1
X_7934_ _3389_ _3448_ _3462_ _3564_ VGND VGND 
+ VPWR
+ VPWR _3565_ sky130_fd_sc_hd__a31o_1
X_7935_ _3460_ _3565_ VGND VGND VPWR VPWR 
+ _3566_
+ sky130_fd_sc_hd__or2_1
X_7936_ _3458_ _3566_ VGND VGND VPWR VPWR 
+ _3567_
+ sky130_fd_sc_hd__or2_1
X_7937_ _3389_ _3448_ _3451_ _3453_ _3567_ VGND 
+ VGND
+ VPWR VPWR _3568_ sky130_fd_sc_hd__a311oi_1
X_7938_ _3447_ _3568_ VGND VGND VPWR VPWR 
+ _3569_
+ sky130_fd_sc_hd__nand2_1
X_7939_ _3442_ _3395_ _3569_ VGND VGND VPWR 
+ VPWR
+ _3570_ sky130_fd_sc_hd__o21ba_1
X_7940_ _3442_ _3444_ _3570_ VGND VGND VPWR 
+ VPWR
+ _3571_ sky130_fd_sc_hd__o21ai_1
X_7941_ _3439_ _3571_ VGND VGND VPWR VPWR 
+ _3572_
+ sky130_fd_sc_hd__or2_1
X_7942_ _3429_ _3434_ _3572_ VGND VGND VPWR 
+ VPWR
+ _3573_ sky130_fd_sc_hd__or3_1
X_7943_ _3392_ _3573_ VGND VGND VPWR VPWR 
+ _3574_
+ sky130_fd_sc_hd__or2_1
X_7944_ _3574_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_7945_ _3478_ _3428_ \wbbd_state[9]\ VGND VGND VPWR 
+ VPWR
+ _3575_ sky130_fd_sc_hd__o21ai_1
X_7946_ _3430_ _3470_ VGND VGND VPWR VPWR 
+ _3576_
+ sky130_fd_sc_hd__or2_1
X_7947_ net156 net153 _3576_ VGND VGND VPWR 
+ VPWR
+ _3577_ sky130_fd_sc_hd__or3_1
X_7948_ _3577_ VGND VGND VPWR VPWR _3578_ sky130_fd_sc_hd__buf_12
X_7949_ _3428_ _3578_ VGND VGND VPWR VPWR 
+ _3579_
+ sky130_fd_sc_hd__or2_1
X_7950_ _3390_ _3472_ _3388_ VGND VGND VPWR 
+ VPWR
+ _3580_ sky130_fd_sc_hd__or3_1
X_7951_ net158 _3424_ _3421_ _3415_ VGND VGND 
+ VPWR
+ VPWR _3581_ sky130_fd_sc_hd__or4_1
X_7952_ _3581_ VGND VGND VPWR VPWR _3582_ sky130_fd_sc_hd__clkbuf_4
X_7953_ _3470_ _3435_ VGND VGND VPWR VPWR 
+ _3583_
+ sky130_fd_sc_hd__or2_1
X_7954_ _3583_ VGND VGND VPWR VPWR _3584_ sky130_fd_sc_hd__buf_12
X_7955_ _3582_ _3584_ VGND VGND VPWR VPWR 
+ _3585_
+ sky130_fd_sc_hd__nor2_2
X_7956_ _3430_ _3393_ _3383_ VGND VGND VPWR 
+ VPWR
+ _3586_ sky130_fd_sc_hd__or3_1
X_7957_ _3404_ _3396_ _3586_ VGND VGND VPWR 
+ VPWR
+ _3587_ sky130_fd_sc_hd__or3_1
X_7958_ _3396_ _3586_ VGND VGND VPWR VPWR 
+ _3588_
+ sky130_fd_sc_hd__or2_1
X_7959_ _3403_ _3404_ _3588_ VGND VGND VPWR 
+ VPWR
+ _3589_ sky130_fd_sc_hd__or3_2
X_7960_ _3589_ VGND VGND VPWR VPWR _3590_ sky130_fd_sc_hd__inv_2
X_7961_ _3403_ _3587_ _3590_ VGND VGND VPWR 
+ VPWR
+ _3591_ sky130_fd_sc_hd__a21oi_1
X_7962_ net160 _3590_ _3400_ _3589_ VGND VGND 
+ VPWR
+ VPWR _3592_ sky130_fd_sc_hd__o22a_1
X_7963_ _3591_ _3592_ VGND VGND VPWR VPWR 
+ _3593_
+ sky130_fd_sc_hd__or2_4
X_7964_ _3396_ _3586_ _3588_ VGND VGND VPWR 
+ VPWR
+ _3594_ sky130_fd_sc_hd__a21bo_2
X_7965_ _3404_ _3594_ VGND VGND VPWR VPWR 
+ _3595_
+ sky130_fd_sc_hd__or2_2
X_7966_ _3399_ _3588_ _3406_ VGND VGND VPWR 
+ VPWR
+ _3596_ sky130_fd_sc_hd__or3_1
X_7967_ _1795_ _3596_ _1795_ _3596_ VGND VGND 
+ VPWR
+ VPWR _3597_ sky130_fd_sc_hd__o2bb2a_1
X_7968_ _3597_ _3413_ VGND VGND VPWR VPWR 
+ _3598_
+ sky130_fd_sc_hd__or2_1
X_7969_ _3411_ _3598_ VGND VGND VPWR VPWR 
+ _3599_
+ sky130_fd_sc_hd__or2_1
X_7970_ _3599_ VGND VGND VPWR VPWR _3600_ sky130_fd_sc_hd__buf_6
X_7971_ _3595_ _3600_ VGND VGND VPWR VPWR 
+ _3601_
+ sky130_fd_sc_hd__or2_1
X_7972_ _3593_ _3601_ VGND VGND VPWR VPWR 
+ _3602_
+ sky130_fd_sc_hd__or2_1
X_7973_ _3602_ VGND VGND VPWR VPWR _3603_ sky130_fd_sc_hd__clkbuf_4
X_7974_ net153 _3431_ VGND VGND VPWR VPWR 
+ _3604_
+ sky130_fd_sc_hd__or2_1
X_7975_ _3604_ VGND VGND VPWR VPWR _3605_ sky130_fd_sc_hd__buf_8
X_7976_ _3404_ _3588_ _3587_ VGND VGND VPWR 
+ VPWR
+ _3606_ sky130_fd_sc_hd__a21bo_1
X_7977_ _3594_ _3606_ VGND VGND VPWR VPWR 
+ _3607_
+ sky130_fd_sc_hd__nand2_4
X_7978_ _3607_ _3600_ VGND VGND VPWR VPWR 
+ _3608_
+ sky130_fd_sc_hd__or2_1
X_7979_ _3591_ VGND VGND VPWR VPWR _3609_ sky130_fd_sc_hd__inv_2
X_7980_ net160 _3609_ VGND VGND VPWR VPWR 
+ _3610_
+ sky130_fd_sc_hd__or2_4
X_7981_ _3608_ _3610_ VGND VGND VPWR VPWR 
+ _3611_
+ sky130_fd_sc_hd__or2_1
X_7982_ _3611_ VGND VGND VPWR VPWR _3612_ sky130_fd_sc_hd__clkbuf_4
X_7983_ _3446_ VGND VGND VPWR VPWR _3613_ sky130_fd_sc_hd__clkinv_4
X_7984_ net158 _3594_ _3600_ VGND VGND VPWR 
+ VPWR
+ _3614_ sky130_fd_sc_hd__or3_2
X_7985_ _3614_ _3610_ VGND VGND VPWR VPWR 
+ _3615_
+ sky130_fd_sc_hd__or2_1
X_7986_ _3615_ VGND VGND VPWR VPWR _3616_ sky130_fd_sc_hd__buf_2
X_7987_ _3616_ VGND VGND VPWR VPWR _3617_ sky130_fd_sc_hd__inv_2
X_7988_ _3606_ _3594_ VGND VGND VPWR VPWR 
+ _3618_
+ sky130_fd_sc_hd__or2b_2
X_7989_ _3600_ _3618_ VGND VGND VPWR VPWR 
+ _3619_
+ sky130_fd_sc_hd__or2_1
X_7990_ _3619_ _3610_ VGND VGND VPWR VPWR 
+ _3620_
+ sky130_fd_sc_hd__or2_1
X_7991_ _3620_ VGND VGND VPWR VPWR _3621_ sky130_fd_sc_hd__clkbuf_4
X_7992_ _3601_ _3610_ VGND VGND VPWR VPWR 
+ _3622_
+ sky130_fd_sc_hd__or2_1
X_7993_ _3622_ VGND VGND VPWR VPWR _3623_ sky130_fd_sc_hd__buf_4
X_7994_ _3609_ _3592_ VGND VGND VPWR VPWR 
+ _3624_
+ sky130_fd_sc_hd__nand2_4
X_7995_ _3624_ _3608_ VGND VGND VPWR VPWR 
+ _3625_
+ sky130_fd_sc_hd__or2_1
X_7996_ _3625_ VGND VGND VPWR VPWR _3626_ sky130_fd_sc_hd__clkbuf_4
X_7997_ _3624_ _3614_ VGND VGND VPWR VPWR 
+ _3627_
+ sky130_fd_sc_hd__or2_1
X_7998_ _3627_ VGND VGND VPWR VPWR _3628_ sky130_fd_sc_hd__clkbuf_4
X_7999_ _3624_ _3619_ VGND VGND VPWR VPWR 
+ _3629_
+ sky130_fd_sc_hd__or2_1
X_8000_ _3629_ VGND VGND VPWR VPWR _3630_ sky130_fd_sc_hd__buf_6
X_8001_ _3446_ _3630_ VGND VGND VPWR VPWR 
+ _3631_
+ sky130_fd_sc_hd__nor2_1
X_8002_ _3390_ _3478_ VGND VGND VPWR VPWR 
+ _3632_
+ sky130_fd_sc_hd__or2_1
X_8003_ _3632_ VGND VGND VPWR VPWR _3633_ sky130_fd_sc_hd__inv_2
X_8004_ _3390_ _3584_ VGND VGND VPWR VPWR 
+ _3634_
+ sky130_fd_sc_hd__or2_1
X_8005_ _3634_ VGND VGND VPWR VPWR _3635_ sky130_fd_sc_hd__inv_2
X_8006_ _3529_ VGND VGND VPWR VPWR _3636_ sky130_fd_sc_hd__clkinv_2
X_8007_ _3633_ _3635_ _3636_ VGND VGND VPWR 
+ VPWR
+ _3637_ sky130_fd_sc_hd__o21a_1
X_8008_ _3413_ _3410_ _3528_ VGND VGND VPWR 
+ VPWR
+ _3638_ sky130_fd_sc_hd__or3_4
X_8009_ _3632_ _3638_ VGND VGND VPWR VPWR 
+ _3639_
+ sky130_fd_sc_hd__or2_1
X_8010_ _3495_ _3426_ _3639_ VGND VGND VPWR 
+ VPWR
+ _3640_ sky130_fd_sc_hd__o21ai_1
X_8011_ _3404_ _3424_ _3529_ VGND VGND VPWR 
+ VPWR
+ _3641_ sky130_fd_sc_hd__or3_2
X_8012_ _3641_ _3531_ VGND VGND VPWR VPWR 
+ _3642_
+ sky130_fd_sc_hd__or2_1
X_8013_ _3446_ _3642_ VGND VGND VPWR VPWR 
+ _3643_
+ sky130_fd_sc_hd__or2_1
X_8014_ _3437_ _3630_ _3643_ VGND VGND VPWR 
+ VPWR
+ _3644_ sky130_fd_sc_hd__o21ai_1
X_8015_ _3532_ _3642_ _3431_ VGND VGND VPWR 
+ VPWR
+ _3645_ sky130_fd_sc_hd__a21oi_1
X_8016_ _3637_ _3640_ _3644_ _3645_ VGND VGND 
+ VPWR
+ VPWR _3646_ sky130_fd_sc_hd__or4_1
X_8017_ _3437_ _3628_ VGND VGND VPWR VPWR 
+ _3647_
+ sky130_fd_sc_hd__or2_1
X_8018_ _3433_ _3628_ VGND VGND VPWR VPWR 
+ _3648_
+ sky130_fd_sc_hd__or2_1
X_8019_ _3631_ _3646_ _3647_ _3648_ VGND VGND 
+ VPWR
+ VPWR _3649_ sky130_fd_sc_hd__and4bb_1
X_8020_ _3628_ _3605_ _3446_ _3628_ _3649_ VGND 
+ VGND
+ VPWR VPWR _3650_ sky130_fd_sc_hd__o221a_1
X_8021_ _3437_ _3626_ VGND VGND VPWR VPWR 
+ _3651_
+ sky130_fd_sc_hd__or2_1
X_8022_ _3433_ _3626_ VGND VGND VPWR VPWR 
+ _3652_
+ sky130_fd_sc_hd__or2_1
X_8023_ _3605_ _3626_ _3650_ _3651_ _3652_ VGND 
+ VGND
+ VPWR VPWR _3653_ sky130_fd_sc_hd__o2111a_1
X_8024_ _3437_ _3623_ VGND VGND VPWR VPWR 
+ _3654_
+ sky130_fd_sc_hd__or2_1
X_8025_ _3433_ _3623_ VGND VGND VPWR VPWR 
+ _3655_
+ sky130_fd_sc_hd__or2_1
X_8026_ _3446_ _3626_ _3653_ _3654_ _3655_ VGND 
+ VGND
+ VPWR VPWR _3656_ sky130_fd_sc_hd__o2111a_1
X_8027_ _3605_ _3623_ _3446_ _3623_ _3656_ VGND 
+ VGND
+ VPWR VPWR _3657_ sky130_fd_sc_hd__o221a_1
X_8028_ _3437_ _3621_ VGND VGND VPWR VPWR 
+ _3658_
+ sky130_fd_sc_hd__or2_1
X_8029_ _3433_ _3621_ VGND VGND VPWR VPWR 
+ _3659_
+ sky130_fd_sc_hd__or2_1
X_8030_ _3605_ _3621_ _3657_ _3658_ _3659_ VGND 
+ VGND
+ VPWR VPWR _3660_ sky130_fd_sc_hd__o2111a_1
X_8031_ _3446_ _3621_ _3660_ VGND VGND VPWR 
+ VPWR
+ _3661_ sky130_fd_sc_hd__o21ai_1
X_8032_ _3437_ _3616_ VGND VGND VPWR VPWR 
+ _3662_
+ sky130_fd_sc_hd__nor2_1
X_8033_ _3661_ _3662_ VGND VGND VPWR VPWR 
+ _3663_
+ sky130_fd_sc_hd__nor2_1
X_8034_ _3433_ _3616_ VGND VGND VPWR VPWR 
+ _3664_
+ sky130_fd_sc_hd__or2_1
X_8035_ _3663_ _3664_ VGND VGND VPWR VPWR 
+ _3665_
+ sky130_fd_sc_hd__and2_1
X_8036_ _3605_ _3616_ _3665_ VGND VGND VPWR 
+ VPWR
+ _3666_ sky130_fd_sc_hd__o21ai_1
X_8037_ _3613_ _3617_ _3666_ VGND VGND VPWR 
+ VPWR
+ _3667_ sky130_fd_sc_hd__a21oi_1
X_8038_ _3437_ _3612_ VGND VGND VPWR VPWR 
+ _3668_
+ sky130_fd_sc_hd__or2_1
X_8039_ _3667_ _3668_ VGND VGND VPWR VPWR 
+ _3669_
+ sky130_fd_sc_hd__nand2_1
X_8040_ _3433_ _3612_ VGND VGND VPWR VPWR 
+ _3670_
+ sky130_fd_sc_hd__nor2_1
X_8041_ _3669_ _3670_ VGND VGND VPWR VPWR 
+ _3671_
+ sky130_fd_sc_hd__nor2_1
X_8042_ _3605_ _3612_ _3671_ VGND VGND VPWR 
+ VPWR
+ _3672_ sky130_fd_sc_hd__o21a_1
X_8043_ _3446_ _3612_ _3672_ VGND VGND VPWR 
+ VPWR
+ _3673_ sky130_fd_sc_hd__o21ai_1
X_8044_ _3437_ _3603_ VGND VGND VPWR VPWR 
+ _3674_
+ sky130_fd_sc_hd__nor2_1
X_8045_ _3673_ _3674_ VGND VGND VPWR VPWR 
+ _3675_
+ sky130_fd_sc_hd__nor2_1
X_8046_ _3433_ _3603_ VGND VGND VPWR VPWR 
+ _3676_
+ sky130_fd_sc_hd__or2_1
X_8047_ _3675_ _3676_ VGND VGND VPWR VPWR 
+ _3677_
+ sky130_fd_sc_hd__and2_1
X_8048_ _3603_ _3605_ _3677_ VGND VGND VPWR 
+ VPWR
+ _3678_ sky130_fd_sc_hd__o21ai_2
X_8049_ _3446_ _3603_ _3678_ VGND VGND VPWR 
+ VPWR
+ _3679_ sky130_fd_sc_hd__o21ba_1
X_8050_ _3593_ _3619_ VGND VGND VPWR VPWR 
+ _3680_
+ sky130_fd_sc_hd__or2_1
X_8051_ _3680_ VGND VGND VPWR VPWR _3681_ sky130_fd_sc_hd__buf_2
X_8052_ _3437_ _3681_ VGND VGND VPWR VPWR 
+ _3682_
+ sky130_fd_sc_hd__or2_1
X_8053_ _3679_ _3682_ VGND VGND VPWR VPWR 
+ _3683_
+ sky130_fd_sc_hd__nand2_1
X_8054_ _3433_ _3681_ VGND VGND VPWR VPWR 
+ _3684_
+ sky130_fd_sc_hd__nor2_1
X_8055_ _3683_ _3684_ VGND VGND VPWR VPWR 
+ _3685_
+ sky130_fd_sc_hd__nor2_1
X_8056_ _3605_ _3681_ VGND VGND VPWR VPWR 
+ _3686_
+ sky130_fd_sc_hd__or2_1
X_8057_ _3685_ _3686_ VGND VGND VPWR VPWR 
+ _3687_
+ sky130_fd_sc_hd__nand2_1
X_8058_ _3481_ VGND VGND VPWR VPWR _3688_ sky130_fd_sc_hd__inv_2
X_8059_ _3426_ VGND VGND VPWR VPWR _3689_ sky130_fd_sc_hd__inv_2
X_8060_ _3638_ VGND VGND VPWR VPWR _3690_ sky130_fd_sc_hd__inv_2
X_8061_ _3688_ _3689_ _3690_ VGND VGND VPWR 
+ VPWR
+ _3691_ sky130_fd_sc_hd__and3_1
X_8062_ _3687_ _3691_ VGND VGND VPWR VPWR 
+ _3692_
+ sky130_fd_sc_hd__or2_1
X_8063_ _3478_ VGND VGND VPWR VPWR _3693_ sky130_fd_sc_hd__clkinv_4
X_8064_ _3693_ _3689_ _3636_ VGND VGND VPWR 
+ VPWR
+ _3694_ sky130_fd_sc_hd__and3_1
X_8065_ _3692_ _3694_ VGND VGND VPWR VPWR 
+ _3695_
+ sky130_fd_sc_hd__or2_1
X_8066_ _3451_ _3693_ _3389_ VGND VGND VPWR 
+ VPWR
+ _3696_ sky130_fd_sc_hd__and3_1
X_8067_ _3695_ _3696_ VGND VGND VPWR VPWR 
+ _3697_
+ sky130_fd_sc_hd__nor2_1
X_8068_ _3456_ _3584_ VGND VGND VPWR VPWR 
+ _3698_
+ sky130_fd_sc_hd__or2_1
X_8069_ _3697_ _3698_ VGND VGND VPWR VPWR 
+ _3699_
+ sky130_fd_sc_hd__nand2_1
X_8070_ _3456_ _3476_ _3699_ VGND VGND VPWR 
+ VPWR
+ _3700_ sky130_fd_sc_hd__o21bai_1
X_8071_ _3442_ _3478_ VGND VGND VPWR VPWR 
+ _3701_
+ sky130_fd_sc_hd__nor2_4
X_8072_ _3476_ _3582_ VGND VGND VPWR VPWR 
+ _3702_
+ sky130_fd_sc_hd__nor2_1
X_8073_ _3701_ _3702_ VGND VGND VPWR VPWR 
+ _3703_
+ sky130_fd_sc_hd__or2_1
X_8074_ _3700_ _3703_ VGND VGND VPWR VPWR 
+ _3704_
+ sky130_fd_sc_hd__or2_1
X_8075_ _3585_ _3704_ VGND VGND VPWR VPWR 
+ _3705_
+ sky130_fd_sc_hd__nor2_1
X_8076_ _3472_ _3582_ _3705_ VGND VGND VPWR 
+ VPWR
+ _3706_ sky130_fd_sc_hd__o21ai_1
X_8077_ _3478_ _3582_ VGND VGND VPWR VPWR 
+ _3707_
+ sky130_fd_sc_hd__nor2_1
X_8078_ _3706_ _3707_ VGND VGND VPWR VPWR 
+ _3708_
+ sky130_fd_sc_hd__nor2_1
X_8079_ net156 _3383_ _3576_ VGND VGND VPWR 
+ VPWR
+ _3709_ sky130_fd_sc_hd__or3_1
X_8080_ _3709_ VGND VGND VPWR VPWR _3710_ sky130_fd_sc_hd__buf_8
X_8081_ _3428_ _3710_ VGND VGND VPWR VPWR 
+ _3711_
+ sky130_fd_sc_hd__or2_1
X_8082_ _3708_ _3711_ VGND VGND VPWR VPWR 
+ _3712_
+ sky130_fd_sc_hd__and2_1
X_8083_ _3579_ _3580_ _3712_ VGND VGND VPWR 
+ VPWR
+ _3713_ sky130_fd_sc_hd__and3_1
X_8084_ _3415_ _3481_ VGND VGND VPWR VPWR 
+ _3714_
+ sky130_fd_sc_hd__or2_1
X_8085_ _3426_ _3714_ VGND VGND VPWR VPWR 
+ _3715_
+ sky130_fd_sc_hd__or2_1
X_8086_ _3713_ _3715_ VGND VGND VPWR VPWR 
+ _3716_
+ sky130_fd_sc_hd__nand2_1
X_8087_ _3575_ _3716_ VGND VGND VPWR VPWR 
+ _3717_
+ sky130_fd_sc_hd__or2b_1
X_8088_ _3428_ _3605_ VGND VGND VPWR VPWR 
+ _3718_
+ sky130_fd_sc_hd__nor2_1
X_8089_ _3410_ _1794_ _3596_ VGND VGND VPWR 
+ VPWR
+ _3719_ sky130_fd_sc_hd__mux2_1
X_8090_ _3413_ _3593_ _3597_ _3719_ VGND VGND 
+ VPWR
+ VPWR _3720_ sky130_fd_sc_hd__or4bb_4
X_8091_ net158 _3594_ _3720_ VGND VGND VPWR 
+ VPWR
+ _3721_ sky130_fd_sc_hd__or3_1
X_8092_ _3721_ VGND VGND VPWR VPWR _3722_ sky130_fd_sc_hd__inv_2
X_8093_ _3431_ _3721_ VGND VGND VPWR VPWR 
+ _3723_
+ sky130_fd_sc_hd__nor2_1
X_8094_ _3447_ VGND VGND VPWR VPWR _3724_ sky130_fd_sc_hd__inv_2
X_8095_ _3437_ _3582_ VGND VGND VPWR VPWR 
+ _3725_
+ sky130_fd_sc_hd__nor2_1
X_8096_ _3607_ _3593_ VGND VGND VPWR VPWR 
+ _3726_
+ sky130_fd_sc_hd__or2_1
X_8097_ _3726_ _3446_ VGND VGND VPWR VPWR 
+ _3727_
+ sky130_fd_sc_hd__or2_1
X_8098_ _3600_ _3727_ VGND VGND VPWR VPWR 
+ _3728_
+ sky130_fd_sc_hd__nor2_1
X_8099_ _3470_ _3586_ VGND VGND VPWR VPWR 
+ _3729_
+ sky130_fd_sc_hd__or2_1
X_8100_ _3729_ VGND VGND VPWR VPWR _3730_ sky130_fd_sc_hd__buf_12
X_8101_ _3730_ VGND VGND VPWR VPWR _3731_ sky130_fd_sc_hd__clkinv_2
X_8102_ _3470_ _3596_ VGND VGND VPWR VPWR 
+ _3732_
+ sky130_fd_sc_hd__or2_1
X_8103_ _3732_ VGND VGND VPWR VPWR _3733_ sky130_fd_sc_hd__inv_2
X_8104_ net144 _3732_ _3411_ _3733_ VGND VGND 
+ VPWR
+ VPWR _3734_ sky130_fd_sc_hd__a22o_1
X_8105_ _1795_ _3733_ net143 _3732_ VGND VGND 
+ VPWR
+ VPWR _3735_ sky130_fd_sc_hd__o22a_1
X_8106_ _3735_ VGND VGND VPWR VPWR _3736_ sky130_fd_sc_hd__inv_2
X_8107_ _3413_ _3734_ _3736_ VGND VGND VPWR 
+ VPWR
+ _3737_ sky130_fd_sc_hd__or3_1
X_8108_ _3737_ VGND VGND VPWR VPWR _3738_ sky130_fd_sc_hd__buf_6
X_8109_ _3738_ VGND VGND VPWR VPWR _3739_ sky130_fd_sc_hd__inv_2
X_8110_ _3731_ _3451_ _3739_ VGND VGND VPWR 
+ VPWR
+ _3740_ sky130_fd_sc_hd__and3_2
X_8111_ _3578_ VGND VGND VPWR VPWR _3741_ sky130_fd_sc_hd__clkinv_4
X_8112_ _3710_ VGND VGND VPWR VPWR _3742_ sky130_fd_sc_hd__inv_4
X_8113_ _3628_ _3578_ VGND VGND VPWR VPWR 
+ _3743_
+ sky130_fd_sc_hd__nor2_1
X_8114_ _3584_ VGND VGND VPWR VPWR _3744_ sky130_fd_sc_hd__inv_2
X_8115_ _3628_ VGND VGND VPWR VPWR _3745_ sky130_fd_sc_hd__inv_2
X_8116_ _3601_ _3624_ VGND VGND VPWR VPWR 
+ _3746_
+ sky130_fd_sc_hd__or2_2
X_8117_ _3630_ _3746_ VGND VGND VPWR VPWR 
+ _3747_
+ sky130_fd_sc_hd__nand2_2
X_8118_ _3393_ net153 _3630_ VGND VGND VPWR 
+ VPWR
+ _3748_ sky130_fd_sc_hd__or3b_1
X_8119_ _3438_ VGND VGND VPWR VPWR _3749_ sky130_fd_sc_hd__inv_2
X_8120_ _3719_ _3598_ VGND VGND VPWR VPWR 
+ _3750_
+ sky130_fd_sc_hd__or2_4
X_8121_ _3513_ _3750_ _3600_ VGND VGND VPWR 
+ VPWR
+ _3751_ sky130_fd_sc_hd__o21ai_1
X_8122_ _3514_ _3512_ _3749_ _3751_ VGND VGND 
+ VPWR
+ VPWR _3752_ sky130_fd_sc_hd__o31a_1
X_8123_ net142 net131 _3747_ _3748_ _3752_ VGND 
+ VGND
+ VPWR VPWR _3753_ sky130_fd_sc_hd__a41o_2
X_8124_ _3744_ _3745_ _3745_ _3742_ _3753_ VGND 
+ VGND
+ VPWR VPWR _3754_ sky130_fd_sc_hd__a221o_1
X_8125_ _3730_ _3628_ VGND VGND VPWR VPWR 
+ _3755_
+ sky130_fd_sc_hd__nor2_1
X_8126_ _3584_ _3626_ VGND VGND VPWR VPWR 
+ _3756_
+ sky130_fd_sc_hd__nor2_1
X_8127_ _3743_ _3754_ _3755_ _3756_ VGND VGND 
+ VPWR
+ VPWR _3757_ sky130_fd_sc_hd__or4_1
X_8128_ _3626_ _3710_ VGND VGND VPWR VPWR 
+ _3758_
+ sky130_fd_sc_hd__nor2_1
X_8129_ _3626_ _3578_ VGND VGND VPWR VPWR 
+ _3759_
+ sky130_fd_sc_hd__nor2_1
X_8130_ _3730_ _3626_ VGND VGND VPWR VPWR 
+ _3760_
+ sky130_fd_sc_hd__nor2_1
X_8131_ _3757_ _3758_ _3759_ _3760_ VGND VGND 
+ VPWR
+ VPWR _3761_ sky130_fd_sc_hd__or4_1
X_8132_ _3584_ _3623_ VGND VGND VPWR VPWR 
+ _3762_
+ sky130_fd_sc_hd__or2_1
X_8133_ _3762_ VGND VGND VPWR VPWR _3763_ sky130_fd_sc_hd__inv_2
X_8134_ _3623_ _3710_ VGND VGND VPWR VPWR 
+ _3764_
+ sky130_fd_sc_hd__nor2_1
X_8135_ _3623_ _3578_ VGND VGND VPWR VPWR 
+ _3765_
+ sky130_fd_sc_hd__nor2_1
X_8136_ _3761_ _3763_ _3764_ _3765_ VGND VGND 
+ VPWR
+ VPWR _3766_ sky130_fd_sc_hd__or4_1
X_8137_ _3730_ _3623_ VGND VGND VPWR VPWR 
+ _3767_
+ sky130_fd_sc_hd__nor2_1
X_8138_ _3584_ _3621_ VGND VGND VPWR VPWR 
+ _3768_
+ sky130_fd_sc_hd__nor2_1
X_8139_ _3621_ _3710_ VGND VGND VPWR VPWR 
+ _3769_
+ sky130_fd_sc_hd__nor2_1
X_8140_ _3766_ _3767_ _3768_ _3769_ VGND VGND 
+ VPWR
+ VPWR _3770_ sky130_fd_sc_hd__or4_1
X_8141_ _3621_ _3578_ VGND VGND VPWR VPWR 
+ _3771_
+ sky130_fd_sc_hd__nor2_1
X_8142_ _3730_ _3621_ VGND VGND VPWR VPWR 
+ _3772_
+ sky130_fd_sc_hd__nor2_1
X_8143_ _3584_ _3616_ VGND VGND VPWR VPWR 
+ _3773_
+ sky130_fd_sc_hd__nor2_1
X_8144_ _3770_ _3771_ _3772_ _3773_ VGND VGND 
+ VPWR
+ VPWR _3774_ sky130_fd_sc_hd__or4_1
X_8145_ _3617_ _3742_ _3774_ VGND VGND VPWR 
+ VPWR
+ _3775_ sky130_fd_sc_hd__a21o_1
X_8146_ _3617_ _3741_ _3775_ VGND VGND VPWR 
+ VPWR
+ _3776_ sky130_fd_sc_hd__a21o_1
X_8147_ _3730_ _3616_ VGND VGND VPWR VPWR 
+ _3777_
+ sky130_fd_sc_hd__nor2_1
X_8148_ _3776_ _3777_ VGND VGND VPWR VPWR 
+ _3778_
+ sky130_fd_sc_hd__or2_1
X_8149_ _3584_ _3612_ VGND VGND VPWR VPWR 
+ _3779_
+ sky130_fd_sc_hd__nor2_1
X_8150_ _3778_ _3779_ VGND VGND VPWR VPWR 
+ _3780_
+ sky130_fd_sc_hd__or2_1
X_8151_ _3612_ _3710_ VGND VGND VPWR VPWR 
+ _3781_
+ sky130_fd_sc_hd__nor2_1
X_8152_ _3780_ _3781_ VGND VGND VPWR VPWR 
+ _3782_
+ sky130_fd_sc_hd__or2_1
X_8153_ _3612_ _3578_ VGND VGND VPWR VPWR 
+ _3783_
+ sky130_fd_sc_hd__nor2_1
X_8154_ _3782_ _3783_ VGND VGND VPWR VPWR 
+ _3784_
+ sky130_fd_sc_hd__or2_1
X_8155_ _3730_ _3612_ VGND VGND VPWR VPWR 
+ _3785_
+ sky130_fd_sc_hd__nor2_1
X_8156_ _3784_ _3785_ VGND VGND VPWR VPWR 
+ _3786_
+ sky130_fd_sc_hd__or2_1
X_8157_ _3584_ _3603_ VGND VGND VPWR VPWR 
+ _3787_
+ sky130_fd_sc_hd__nor2_1
X_8158_ _3786_ _3787_ VGND VGND VPWR VPWR 
+ _3788_
+ sky130_fd_sc_hd__or2_1
X_8159_ _3603_ _3710_ VGND VGND VPWR VPWR 
+ _3789_
+ sky130_fd_sc_hd__nor2_1
X_8160_ _3788_ _3789_ VGND VGND VPWR VPWR 
+ _3790_
+ sky130_fd_sc_hd__or2_1
X_8161_ _3603_ _3578_ VGND VGND VPWR VPWR 
+ _3791_
+ sky130_fd_sc_hd__nor2_1
X_8162_ _3790_ _3791_ VGND VGND VPWR VPWR 
+ _3792_
+ sky130_fd_sc_hd__or2_1
X_8163_ _3740_ _3792_ VGND VGND VPWR VPWR 
+ _3793_
+ sky130_fd_sc_hd__or2_1
X_8164_ _3584_ _3681_ VGND VGND VPWR VPWR 
+ _3794_
+ sky130_fd_sc_hd__nor2_1
X_8165_ _3793_ _3794_ VGND VGND VPWR VPWR 
+ _3795_
+ sky130_fd_sc_hd__or2_1
X_8166_ _3681_ _3710_ VGND VGND VPWR VPWR 
+ _3796_
+ sky130_fd_sc_hd__nor2_1
X_8167_ _3795_ _3796_ VGND VGND VPWR VPWR 
+ _3797_
+ sky130_fd_sc_hd__or2_1
X_8168_ _3681_ _3578_ VGND VGND VPWR VPWR 
+ _3798_
+ sky130_fd_sc_hd__or2_1
X_8169_ _3798_ VGND VGND VPWR VPWR _3799_ sky130_fd_sc_hd__inv_2
X_8170_ _3726_ _3605_ VGND VGND VPWR VPWR 
+ _3800_
+ sky130_fd_sc_hd__or2_1
X_8171_ _3800_ _3750_ VGND VGND VPWR VPWR 
+ _3801_
+ sky130_fd_sc_hd__or2_1
X_8172_ _3797_ _3799_ _3801_ VGND VGND VPWR 
+ VPWR
+ _3802_ sky130_fd_sc_hd__or3b_1
X_8173_ _3728_ _3802_ VGND VGND VPWR VPWR 
+ _3803_
+ sky130_fd_sc_hd__or2_1
X_8174_ _3460_ _3803_ VGND VGND VPWR VPWR 
+ _3804_
+ sky130_fd_sc_hd__nor2_1
X_8175_ _3457_ _3804_ VGND VGND VPWR VPWR 
+ _3805_
+ sky130_fd_sc_hd__nand2_1
X_8176_ _3437_ _3456_ _3805_ VGND VGND VPWR 
+ VPWR
+ _3806_ sky130_fd_sc_hd__o21bai_1
X_8177_ _3724_ _3725_ _3806_ VGND VGND VPWR 
+ VPWR
+ _3807_ sky130_fd_sc_hd__or3_1
X_8178_ _3453_ _3807_ VGND VGND VPWR VPWR 
+ _3808_
+ sky130_fd_sc_hd__or2_1
X_8179_ net153 _3723_ _3808_ VGND VGND VPWR 
+ VPWR
+ _3809_ sky130_fd_sc_hd__a21o_1
X_8180_ _3613_ _3722_ _3809_ VGND VGND VPWR 
+ VPWR
+ _3810_ sky130_fd_sc_hd__a21oi_1
X_8181_ _3429_ _3434_ _3392_ _3810_ VGND VGND 
+ VPWR
+ VPWR _3811_ sky130_fd_sc_hd__or4b_1
X_8182_ _3718_ _3811_ VGND VGND VPWR VPWR 
+ _3812_
+ sky130_fd_sc_hd__nor2_1
X_8183_ _3607_ _3720_ _3446_ \wbbd_state[7]\ VGND VGND 
+ VPWR
+ VPWR _3813_ sky130_fd_sc_hd__o31ai_4
X_8184_ _3812_ _3813_ VGND VGND VPWR VPWR 
+ _3814_
+ sky130_fd_sc_hd__or2_1
X_8185_ _3579_ VGND VGND VPWR VPWR _3815_ sky130_fd_sc_hd__inv_2
X_8186_ _3711_ VGND VGND VPWR VPWR _3816_ sky130_fd_sc_hd__clkinv_2
X_8187_ _3580_ VGND VGND VPWR VPWR _3817_ sky130_fd_sc_hd__inv_2
X_8188_ _3476_ _3428_ VGND VGND VPWR VPWR 
+ _3818_
+ sky130_fd_sc_hd__nor2_2
X_8189_ _3396_ _3730_ VGND VGND VPWR VPWR 
+ _3819_
+ sky130_fd_sc_hd__nor2_1
X_8190_ _3396_ _3730_ _3819_ VGND VGND VPWR 
+ VPWR
+ _3820_ sky130_fd_sc_hd__a21oi_1
X_8191_ _3820_ VGND VGND VPWR VPWR _3821_ sky130_fd_sc_hd__inv_2
X_8192_ _3470_ _3589_ _3400_ VGND VGND VPWR 
+ VPWR
+ _3822_ sky130_fd_sc_hd__o21a_1
X_8193_ _3400_ _3589_ _3470_ VGND VGND VPWR 
+ VPWR
+ _3823_ sky130_fd_sc_hd__or3_2
X_8194_ _3823_ VGND VGND VPWR VPWR _3824_ sky130_fd_sc_hd__inv_2
X_8195_ _3470_ _3587_ VGND VGND VPWR VPWR 
+ _3825_
+ sky130_fd_sc_hd__nor2_1
X_8196_ net159 _3825_ net131 _3590_ VGND VGND 
+ VPWR
+ VPWR _3826_ sky130_fd_sc_hd__a2bb2o_1
X_8197_ _3822_ _3824_ _3826_ VGND VGND VPWR 
+ VPWR
+ _3827_ sky130_fd_sc_hd__o21ai_2
X_8198_ net158 _3821_ _3827_ VGND VGND VPWR 
+ VPWR
+ _3828_ sky130_fd_sc_hd__or3_1
X_8199_ _3828_ VGND VGND VPWR VPWR _3829_ sky130_fd_sc_hd__clkinvlp_2
X_8200_ _3413_ _3734_ _3735_ VGND VGND VPWR 
+ VPWR
+ _3830_ sky130_fd_sc_hd__or3_2
X_8201_ _3830_ VGND VGND VPWR VPWR _3831_ sky130_fd_sc_hd__inv_2
X_8202_ _3442_ _3730_ VGND VGND VPWR VPWR 
+ _3832_
+ sky130_fd_sc_hd__nor2_4
X_8203_ _3698_ VGND VGND VPWR VPWR _3833_ sky130_fd_sc_hd__inv_2
X_8204_ _3823_ _3738_ VGND VGND VPWR VPWR 
+ _3834_
+ sky130_fd_sc_hd__nor2_1
X_8205_ _3395_ _3521_ _3464_ VGND VGND VPWR 
+ VPWR
+ _3835_ sky130_fd_sc_hd__nor3_2
X_8206_ _3452_ _3464_ VGND VGND VPWR VPWR 
+ _3836_
+ sky130_fd_sc_hd__or2_1
X_8207_ _3836_ VGND VGND VPWR VPWR _3837_ sky130_fd_sc_hd__buf_6
X_8208_ _3521_ _3837_ VGND VGND VPWR VPWR 
+ _3838_
+ sky130_fd_sc_hd__nor2_1
X_8209_ _3385_ _3464_ VGND VGND VPWR VPWR 
+ _3839_
+ sky130_fd_sc_hd__or2_1
X_8210_ _3839_ VGND VGND VPWR VPWR _3840_ sky130_fd_sc_hd__buf_4
X_8211_ _3526_ _3837_ VGND VGND VPWR VPWR 
+ _3841_
+ sky130_fd_sc_hd__or2_2
X_8212_ _3526_ _3840_ _3841_ VGND VGND VPWR 
+ VPWR
+ _3842_ sky130_fd_sc_hd__o21ai_1
X_8213_ _3730_ _3828_ VGND VGND VPWR VPWR 
+ _3843_
+ sky130_fd_sc_hd__or2_1
X_8214_ _3843_ VGND VGND VPWR VPWR _3844_ sky130_fd_sc_hd__inv_2
X_8215_ _3385_ _3535_ VGND VGND VPWR VPWR 
+ _3845_
+ sky130_fd_sc_hd__or2_2
X_8216_ _3395_ _3526_ VGND VGND VPWR VPWR 
+ _3846_
+ sky130_fd_sc_hd__or2_2
X_8217_ _3444_ _3526_ _3632_ _3845_ _3846_ VGND 
+ VGND
+ VPWR VPWR _3847_ sky130_fd_sc_hd__o2111ai_1
X_8218_ _3413_ _3410_ _3736_ VGND VGND VPWR 
+ VPWR
+ _3848_ sky130_fd_sc_hd__or3_2
X_8219_ _3848_ _3843_ VGND VGND VPWR VPWR 
+ _3849_
+ sky130_fd_sc_hd__nor2_1
X_8220_ _3635_ _3844_ _3847_ _3739_ _3849_ VGND 
+ VGND
+ VPWR VPWR _3850_ sky130_fd_sc_hd__o32a_2
X_8221_ _3395_ _3535_ _3738_ VGND VGND VPWR 
+ VPWR
+ _3851_ sky130_fd_sc_hd__or3_1
X_8222_ _3444_ _3535_ _3738_ VGND VGND VPWR 
+ VPWR
+ _3852_ sky130_fd_sc_hd__or3_1
X_8223_ _3851_ _3852_ VGND VGND VPWR VPWR 
+ _3853_
+ sky130_fd_sc_hd__and2_1
X_8224_ _3838_ _3842_ _3850_ _3853_ VGND VGND 
+ VPWR
+ VPWR _3854_ sky130_fd_sc_hd__or4b_2
X_8225_ _3521_ _3840_ VGND VGND VPWR VPWR 
+ _3855_
+ sky130_fd_sc_hd__nor2_2
X_8226_ _3444_ _3521_ _3464_ VGND VGND VPWR 
+ VPWR
+ _3856_ sky130_fd_sc_hd__nor3_1
X_8227_ _3835_ _3854_ _3855_ _3856_ VGND VGND 
+ VPWR
+ VPWR _3857_ sky130_fd_sc_hd__or4_1
X_8228_ _3506_ _3837_ VGND VGND VPWR VPWR 
+ _3858_
+ sky130_fd_sc_hd__nor2_2
X_8229_ _3395_ _3507_ VGND VGND VPWR VPWR 
+ _3859_
+ sky130_fd_sc_hd__nor2_1
X_8230_ _3506_ _3840_ VGND VGND VPWR VPWR 
+ _3860_
+ sky130_fd_sc_hd__nor2_1
X_8231_ _3857_ _3858_ _3859_ _3860_ VGND VGND 
+ VPWR
+ VPWR _3861_ sky130_fd_sc_hd__or4_1
X_8232_ _3444_ _3507_ VGND VGND VPWR VPWR 
+ _3862_
+ sky130_fd_sc_hd__or2_1
X_8233_ _3862_ VGND VGND VPWR VPWR _3863_ sky130_fd_sc_hd__inv_2
X_8234_ _3504_ _3837_ VGND VGND VPWR VPWR 
+ _3864_
+ sky130_fd_sc_hd__nor2_1
X_8235_ _3395_ _3505_ VGND VGND VPWR VPWR 
+ _3865_
+ sky130_fd_sc_hd__or2_1
X_8236_ _3865_ VGND VGND VPWR VPWR _3866_ sky130_fd_sc_hd__inv_2
X_8237_ _3861_ _3863_ _3864_ _3866_ VGND VGND 
+ VPWR
+ VPWR _3867_ sky130_fd_sc_hd__or4_1
X_8238_ _3504_ _3840_ VGND VGND VPWR VPWR 
+ _3868_
+ sky130_fd_sc_hd__nor2_1
X_8239_ _3444_ _3505_ VGND VGND VPWR VPWR 
+ _3869_
+ sky130_fd_sc_hd__nor2_1
X_8240_ _3499_ _3837_ VGND VGND VPWR VPWR 
+ _3870_
+ sky130_fd_sc_hd__nor2_1
X_8241_ _3867_ _3868_ _3869_ _3870_ VGND VGND 
+ VPWR
+ VPWR _3871_ sky130_fd_sc_hd__or4_1
X_8242_ _3395_ _3501_ VGND VGND VPWR VPWR 
+ _3872_
+ sky130_fd_sc_hd__or2_1
X_8243_ _3872_ VGND VGND VPWR VPWR _3873_ sky130_fd_sc_hd__inv_2
X_8244_ _3499_ _3840_ VGND VGND VPWR VPWR 
+ _3874_
+ sky130_fd_sc_hd__nor2_1
X_8245_ _3871_ _3873_ _3874_ VGND VGND VPWR 
+ VPWR
+ _3875_ sky130_fd_sc_hd__or3_1
X_8246_ _3444_ _3501_ VGND VGND VPWR VPWR 
+ _3876_
+ sky130_fd_sc_hd__nor2_1
X_8247_ _3497_ _3837_ VGND VGND VPWR VPWR 
+ _3877_
+ sky130_fd_sc_hd__nor2_1
X_8248_ _3875_ _3876_ _3877_ VGND VGND VPWR 
+ VPWR
+ _3878_ sky130_fd_sc_hd__or3_1
X_8249_ _3395_ _3546_ VGND VGND VPWR VPWR 
+ _3879_
+ sky130_fd_sc_hd__or2_1
X_8250_ _3879_ VGND VGND VPWR VPWR _3880_ sky130_fd_sc_hd__inv_2
X_8251_ _3878_ _3880_ VGND VGND VPWR VPWR 
+ _3881_
+ sky130_fd_sc_hd__or2_1
X_8252_ _3497_ _3840_ VGND VGND VPWR VPWR 
+ _3882_
+ sky130_fd_sc_hd__nor2_1
X_8253_ _3881_ _3882_ VGND VGND VPWR VPWR 
+ _3883_
+ sky130_fd_sc_hd__or2_1
X_8254_ _3444_ _3546_ VGND VGND VPWR VPWR 
+ _3884_
+ sky130_fd_sc_hd__nor2_1
X_8255_ _3883_ _3884_ VGND VGND VPWR VPWR 
+ _3885_
+ sky130_fd_sc_hd__or2_1
X_8256_ _3487_ _3837_ VGND VGND VPWR VPWR 
+ _3886_
+ sky130_fd_sc_hd__nor2_1
X_8257_ _3885_ _3886_ VGND VGND VPWR VPWR 
+ _3887_
+ sky130_fd_sc_hd__or2_1
X_8258_ _3395_ _3489_ VGND VGND VPWR VPWR 
+ _3888_
+ sky130_fd_sc_hd__nor2_1
X_8259_ _3887_ _3888_ VGND VGND VPWR VPWR 
+ _3889_
+ sky130_fd_sc_hd__or2_1
X_8260_ _3487_ _3840_ VGND VGND VPWR VPWR 
+ _3890_
+ sky130_fd_sc_hd__nor2_1
X_8261_ _3889_ _3890_ VGND VGND VPWR VPWR 
+ _3891_
+ sky130_fd_sc_hd__or2_1
X_8262_ _3444_ _3489_ VGND VGND VPWR VPWR 
+ _3892_
+ sky130_fd_sc_hd__nor2_1
X_8263_ _3891_ _3892_ VGND VGND VPWR VPWR 
+ _3893_
+ sky130_fd_sc_hd__or2_1
X_8264_ _3461_ _3837_ VGND VGND VPWR VPWR 
+ _3894_
+ sky130_fd_sc_hd__nor2_1
X_8265_ _3893_ _3894_ VGND VGND VPWR VPWR 
+ _3895_
+ sky130_fd_sc_hd__or2_1
X_8266_ _3395_ _3483_ VGND VGND VPWR VPWR 
+ _3896_
+ sky130_fd_sc_hd__nor2_1
X_8267_ _3895_ _3896_ VGND VGND VPWR VPWR 
+ _3897_
+ sky130_fd_sc_hd__or2_1
X_8268_ _3385_ _3483_ VGND VGND VPWR VPWR 
+ _3898_
+ sky130_fd_sc_hd__nor2_1
X_8269_ _3897_ _3898_ VGND VGND VPWR VPWR 
+ _3899_
+ sky130_fd_sc_hd__or2_1
X_8270_ _3444_ _3483_ VGND VGND VPWR VPWR 
+ _3900_
+ sky130_fd_sc_hd__nor2_1
X_8271_ _3899_ _3900_ VGND VGND VPWR VPWR 
+ _3901_
+ sky130_fd_sc_hd__or2_1
X_8272_ _3452_ _3450_ _3465_ VGND VGND VPWR 
+ VPWR
+ _3902_ sky130_fd_sc_hd__nor3_1
X_8273_ _3901_ _3902_ VGND VGND VPWR VPWR 
+ _3903_
+ sky130_fd_sc_hd__or2_1
X_8274_ _3395_ _3450_ _3465_ VGND VGND VPWR 
+ VPWR
+ _3904_ sky130_fd_sc_hd__nor3_1
X_8275_ _3903_ _3904_ VGND VGND VPWR VPWR 
+ _3905_
+ sky130_fd_sc_hd__or2_2
X_8276_ _3385_ _3450_ _3465_ VGND VGND VPWR 
+ VPWR
+ _3906_ sky130_fd_sc_hd__or3_2
X_8277_ net158 _3396_ _3730_ _3404_ _3819_ VGND 
+ VGND
+ VPWR VPWR _3907_ sky130_fd_sc_hd__o32a_1
X_8278_ _3820_ _3827_ _3907_ VGND VGND VPWR 
+ VPWR
+ _3908_ sky130_fd_sc_hd__or3b_1
X_8279_ _3908_ _3578_ _3848_ VGND VGND VPWR 
+ VPWR
+ _3909_ sky130_fd_sc_hd__or3_1
X_8280_ _3905_ _3906_ _3909_ VGND VGND VPWR 
+ VPWR
+ _3910_ sky130_fd_sc_hd__nand3b_1
X_8281_ _3834_ _3910_ VGND VGND VPWR VPWR 
+ _3911_
+ sky130_fd_sc_hd__or2_1
X_8282_ _3731_ _3451_ _3389_ VGND VGND VPWR 
+ VPWR
+ _3912_ sky130_fd_sc_hd__and3_1
X_8283_ _3911_ _3912_ VGND VGND VPWR VPWR 
+ _3913_
+ sky130_fd_sc_hd__or2_1
X_8284_ _3696_ _3913_ VGND VGND VPWR VPWR 
+ _3914_
+ sky130_fd_sc_hd__or2_1
X_8285_ _3833_ _3914_ VGND VGND VPWR VPWR 
+ _3915_
+ sky130_fd_sc_hd__or2_1
X_8286_ _3585_ _3832_ _3915_ VGND VGND VPWR 
+ VPWR
+ _3916_ sky130_fd_sc_hd__or3_1
X_8287_ _3701_ _3916_ VGND VGND VPWR VPWR 
+ _3917_
+ sky130_fd_sc_hd__or2_1
X_8288_ _3831_ _3742_ _3829_ _3917_ VGND VGND 
+ VPWR
+ VPWR _3918_ sky130_fd_sc_hd__a31o_1
X_8289_ _3731_ _3829_ _3831_ _3918_ VGND VGND 
+ VPWR
+ VPWR _3919_ sky130_fd_sc_hd__a31o_1
X_8290_ _3818_ _3919_ VGND VGND VPWR VPWR 
+ _3920_
+ sky130_fd_sc_hd__or2_1
X_8291_ _3816_ _3817_ _3920_ VGND VGND VPWR 
+ VPWR
+ _3921_ sky130_fd_sc_hd__or3_1
X_8292_ _3815_ _3921_ VGND VGND VPWR VPWR 
+ _3922_
+ sky130_fd_sc_hd__nor2_1
X_8293_ _3830_ _3823_ \wbbd_state[8]\ VGND VGND VPWR 
+ VPWR
+ _3923_ sky130_fd_sc_hd__o21ai_2
X_8294_ _3922_ _3923_ VGND VGND VPWR VPWR 
+ _3924_
+ sky130_fd_sc_hd__or2_1
X_8295_ _3814_ _3924_ VGND VGND VPWR VPWR 
+ _3925_
+ sky130_fd_sc_hd__and2_1
X_8296_ _3717_ _3925_ VGND VGND VPWR VPWR 
+ _0179_
+ sky130_fd_sc_hd__nand2_1
X_8297_ _3429_ _3818_ VGND VGND VPWR VPWR 
+ _3926_
+ sky130_fd_sc_hd__or2_1
X_8298_ _3469_ VGND VGND VPWR VPWR _3927_ sky130_fd_sc_hd__inv_2
X_8299_ _3386_ _3492_ VGND VGND VPWR VPWR 
+ _3928_
+ sky130_fd_sc_hd__nor2_1
X_8300_ _3465_ _3928_ VGND VGND VPWR VPWR 
+ _3929_
+ sky130_fd_sc_hd__or2_1
X_8301_ _3929_ VGND VGND VPWR VPWR _3930_ sky130_fd_sc_hd__buf_6
X_8302_ _3930_ VGND VGND VPWR VPWR _3931_ sky130_fd_sc_hd__inv_2
X_8303_ _3539_ VGND VGND VPWR VPWR _3932_ sky130_fd_sc_hd__inv_2
X_8304_ _3932_ _3864_ VGND VGND VPWR VPWR 
+ _3933_
+ sky130_fd_sc_hd__nor2_1
X_8305_ _3476_ _3521_ VGND VGND VPWR VPWR 
+ _3934_
+ sky130_fd_sc_hd__or2_1
X_8306_ _3481_ _3515_ _3934_ _3845_ _3513_ VGND 
+ VGND
+ VPWR VPWR _3935_ sky130_fd_sc_hd__o2111a_1
X_8307_ _3521_ _3837_ _3522_ VGND VGND VPWR 
+ VPWR
+ _3936_ sky130_fd_sc_hd__o21ai_1
X_8308_ _3391_ _3386_ _3466_ _3510_ VGND VGND 
+ VPWR
+ VPWR _3937_ sky130_fd_sc_hd__a31o_1
X_8309_ _3495_ _3535_ _3526_ _3930_ VGND VGND 
+ VPWR
+ VPWR _3938_ sky130_fd_sc_hd__o22a_1
X_8310_ _3855_ _3936_ _3937_ _3938_ VGND VGND 
+ VPWR
+ VPWR _3939_ sky130_fd_sc_hd__or4b_1
X_8311_ _3738_ _3843_ VGND VGND VPWR VPWR 
+ _3940_
+ sky130_fd_sc_hd__or2_2
X_8312_ _3939_ _3858_ _3940_ _3841_ VGND VGND 
+ VPWR
+ VPWR _3941_ sky130_fd_sc_hd__and4bb_1
X_8313_ _3465_ _3935_ _3506_ _3930_ _3941_ VGND 
+ VGND
+ VPWR VPWR _3942_ sky130_fd_sc_hd__o221a_2
X_8314_ _3499_ _3837_ _3542_ VGND VGND VPWR 
+ VPWR
+ _3943_ sky130_fd_sc_hd__o21a_1
X_8315_ _3504_ _3930_ _3933_ _3942_ _3943_ VGND 
+ VGND
+ VPWR VPWR _3944_ sky130_fd_sc_hd__o2111ai_1
X_8316_ _3499_ _3930_ VGND VGND VPWR VPWR 
+ _3945_
+ sky130_fd_sc_hd__nor2_1
X_8317_ _3545_ _3877_ VGND VGND VPWR VPWR 
+ _3946_
+ sky130_fd_sc_hd__or2_1
X_8318_ _3944_ _3945_ _3946_ VGND VGND VPWR 
+ VPWR
+ _3947_ sky130_fd_sc_hd__or3_1
X_8319_ _3497_ _3930_ VGND VGND VPWR VPWR 
+ _3948_
+ sky130_fd_sc_hd__nor2_1
X_8320_ _3550_ VGND VGND VPWR VPWR _3949_ sky130_fd_sc_hd__inv_2
X_8321_ _3949_ _3886_ VGND VGND VPWR VPWR 
+ _3950_
+ sky130_fd_sc_hd__or2_1
X_8322_ _3493_ _3931_ _3947_ _3948_ _3950_ VGND 
+ VGND
+ VPWR VPWR _3951_ sky130_fd_sc_hd__a2111o_2
X_8323_ _3490_ _3894_ VGND VGND VPWR VPWR 
+ _3952_
+ sky130_fd_sc_hd__or2_1
X_8324_ _3461_ _3930_ VGND VGND VPWR VPWR 
+ _3953_
+ sky130_fd_sc_hd__nor2_1
X_8325_ _3484_ VGND VGND VPWR VPWR _3954_ sky130_fd_sc_hd__inv_2
X_8326_ _3954_ _3902_ VGND VGND VPWR VPWR 
+ _3955_
+ sky130_fd_sc_hd__or2_1
X_8327_ _3951_ _3952_ _3953_ _3955_ VGND VGND 
+ VPWR
+ VPWR _3956_ sky130_fd_sc_hd__nor4_2
X_8328_ _3473_ _3928_ _3956_ VGND VGND VPWR 
+ VPWR
+ _3957_ sky130_fd_sc_hd__o21ai_1
X_8329_ _3467_ _3927_ _3957_ VGND VGND VPWR 
+ VPWR
+ _3958_ sky130_fd_sc_hd__or3_1
X_8330_ _3460_ _3912_ VGND VGND VPWR VPWR 
+ _3959_
+ sky130_fd_sc_hd__or2_1
X_8331_ _3958_ _3959_ VGND VGND VPWR VPWR 
+ _3960_
+ sky130_fd_sc_hd__or2_1
X_8332_ _3386_ _3389_ _3451_ _3960_ VGND VGND 
+ VPWR
+ VPWR _3961_ sky130_fd_sc_hd__a31o_1
X_8333_ _3724_ _3701_ _3961_ VGND VGND VPWR 
+ VPWR
+ _3962_ sky130_fd_sc_hd__or3_1
X_8334_ _3442_ _3395_ _3385_ _3442_ VGND VGND 
+ VPWR
+ VPWR _3963_ sky130_fd_sc_hd__o22a_1
X_8335_ _3962_ _3963_ VGND VGND VPWR VPWR 
+ _3964_
+ sky130_fd_sc_hd__or2b_1
X_8336_ _3926_ _3964_ VGND VGND VPWR VPWR 
+ _3965_
+ sky130_fd_sc_hd__or2_1
X_8337_ _3392_ _3817_ _3965_ VGND VGND VPWR 
+ VPWR
+ _3966_ sky130_fd_sc_hd__or3_1
X_8338_ _3966_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
X_8339_ _3429_ _3816_ VGND VGND VPWR VPWR 
+ _3967_
+ sky130_fd_sc_hd__or2_2
X_8340_ _3576_ _3829_ _3831_ _3393_ VGND VGND 
+ VPWR
+ VPWR _3968_ sky130_fd_sc_hd__and4b_1
X_8341_ _3444_ _3526_ _3465_ VGND VGND VPWR 
+ VPWR
+ _3969_ sky130_fd_sc_hd__nor3_1
X_8342_ _3744_ _3745_ _3969_ VGND VGND VPWR 
+ VPWR
+ _3970_ sky130_fd_sc_hd__a21o_1
X_8343_ _3514_ _3633_ _3739_ VGND VGND VPWR 
+ VPWR
+ _3971_ sky130_fd_sc_hd__o21ai_2
X_8344_ _3908_ _3578_ _3738_ _3848_ _3843_ VGND 
+ VGND
+ VPWR VPWR _3972_ sky130_fd_sc_hd__o32a_2
X_8345_ _3820_ _3907_ VGND VGND VPWR VPWR 
+ _3973_
+ sky130_fd_sc_hd__or2_1
X_8346_ _3822_ _3824_ _3826_ VGND VGND VPWR 
+ VPWR
+ _3974_ sky130_fd_sc_hd__or3b_1
X_8347_ _3973_ _3974_ VGND VGND VPWR VPWR 
+ _3975_
+ sky130_fd_sc_hd__or2_2
X_8348_ _3578_ _3975_ _3846_ VGND VGND VPWR 
+ VPWR
+ _3976_ sky130_fd_sc_hd__o21a_1
X_8349_ _3738_ _3976_ VGND VGND VPWR VPWR 
+ _3977_
+ sky130_fd_sc_hd__or2_2
X_8350_ _3404_ _3821_ _3974_ VGND VGND VPWR 
+ VPWR
+ _3978_ sky130_fd_sc_hd__or3_4
X_8351_ _3738_ _3578_ _3978_ VGND VGND VPWR 
+ VPWR
+ _3979_ sky130_fd_sc_hd__or3_1
X_8352_ _3972_ _3977_ _3979_ VGND VGND VPWR 
+ VPWR
+ _3980_ sky130_fd_sc_hd__and3_1
X_8353_ _3584_ _3630_ _3971_ _3853_ _3980_ VGND 
+ VGND
+ VPWR VPWR _3981_ sky130_fd_sc_hd__o2111ai_4
X_8354_ _3743_ _3835_ VGND VGND VPWR VPWR 
+ _3982_
+ sky130_fd_sc_hd__or2_1
X_8355_ _3756_ _3856_ VGND VGND VPWR VPWR 
+ _3983_
+ sky130_fd_sc_hd__or2_1
X_8356_ _3970_ _3981_ _3982_ _3983_ VGND VGND 
+ VPWR
+ VPWR _3984_ sky130_fd_sc_hd__or4_1
X_8357_ _3759_ _3859_ VGND VGND VPWR VPWR 
+ _3985_
+ sky130_fd_sc_hd__or2_1
X_8358_ _3763_ _3863_ VGND VGND VPWR VPWR 
+ _3986_
+ sky130_fd_sc_hd__or2_1
X_8359_ _3765_ _3866_ VGND VGND VPWR VPWR 
+ _3987_
+ sky130_fd_sc_hd__or2_1
X_8360_ _3984_ _3985_ _3986_ _3987_ VGND VGND 
+ VPWR
+ VPWR _3988_ sky130_fd_sc_hd__or4_1
X_8361_ _3768_ _3869_ VGND VGND VPWR VPWR 
+ _3989_
+ sky130_fd_sc_hd__or2_1
X_8362_ _3771_ _3873_ VGND VGND VPWR VPWR 
+ _3990_
+ sky130_fd_sc_hd__or2_1
X_8363_ _3773_ _3876_ VGND VGND VPWR VPWR 
+ _3991_
+ sky130_fd_sc_hd__or2_1
X_8364_ _3988_ _3989_ _3990_ _3991_ VGND VGND 
+ VPWR
+ VPWR _3992_ sky130_fd_sc_hd__or4_1
X_8365_ _3616_ _3578_ _3879_ VGND VGND VPWR 
+ VPWR
+ _3993_ sky130_fd_sc_hd__o21ai_1
X_8366_ _3779_ _3884_ VGND VGND VPWR VPWR 
+ _3994_
+ sky130_fd_sc_hd__or2_1
X_8367_ _3783_ _3888_ VGND VGND VPWR VPWR 
+ _3995_
+ sky130_fd_sc_hd__or2_1
X_8368_ _3992_ _3993_ _3994_ _3995_ VGND VGND 
+ VPWR
+ VPWR _3996_ sky130_fd_sc_hd__or4_2
X_8369_ _3787_ _3892_ VGND VGND VPWR VPWR 
+ _3997_
+ sky130_fd_sc_hd__or2_1
X_8370_ _3791_ _3896_ VGND VGND VPWR VPWR 
+ _3998_
+ sky130_fd_sc_hd__or2_1
X_8371_ _3794_ _3900_ VGND VGND VPWR VPWR 
+ _3999_
+ sky130_fd_sc_hd__or2_1
X_8372_ _3996_ _3997_ _3998_ _3999_ VGND VGND 
+ VPWR
+ VPWR _4000_ sky130_fd_sc_hd__or4_4
X_8373_ _3799_ _3904_ VGND VGND VPWR VPWR 
+ _4001_
+ sky130_fd_sc_hd__or2_2
X_8374_ _3823_ _3848_ _3909_ VGND VGND VPWR 
+ VPWR
+ _4002_ sky130_fd_sc_hd__o21ai_1
X_8375_ _4000_ _4001_ _3834_ _4002_ VGND VGND 
+ VPWR
+ VPWR _4003_ sky130_fd_sc_hd__or4_1
X_8376_ _3460_ _3696_ VGND VGND VPWR VPWR 
+ _4004_
+ sky130_fd_sc_hd__or2_1
X_8377_ _3827_ _3973_ _3830_ VGND VGND VPWR 
+ VPWR
+ _4005_ sky130_fd_sc_hd__or3_1
X_8378_ _4005_ _3578_ VGND VGND VPWR VPWR 
+ _4006_
+ sky130_fd_sc_hd__nor2_1
X_8379_ _3442_ net153 _3430_ net156 VGND VGND 
+ VPWR
+ VPWR _4007_ sky130_fd_sc_hd__and4b_1
X_8380_ _4003_ _4004_ _4006_ _4007_ VGND VGND 
+ VPWR
+ VPWR _4008_ sky130_fd_sc_hd__or4_1
X_8381_ _3968_ _4008_ VGND VGND VPWR VPWR 
+ _4009_
+ sky130_fd_sc_hd__or2_1
X_8382_ _3967_ _4009_ VGND VGND VPWR VPWR 
+ _4010_
+ sky130_fd_sc_hd__or2_1
X_8383_ _3392_ _3815_ VGND VGND VPWR VPWR 
+ _4011_
+ sky130_fd_sc_hd__or2_1
X_8384_ _4010_ _4011_ VGND VGND VPWR VPWR 
+ _4012_
+ sky130_fd_sc_hd__nor2_1
X_8385_ _3923_ _4012_ VGND VGND VPWR VPWR 
+ _4013_
+ sky130_fd_sc_hd__or2_1
X_8386_ _3720_ _3618_ VGND VGND VPWR VPWR 
+ _4014_
+ sky130_fd_sc_hd__or2_1
X_8387_ _3605_ _4014_ VGND VGND VPWR VPWR 
+ _4015_
+ sky130_fd_sc_hd__nor2_1
X_8388_ _3727_ _3750_ _3801_ VGND VGND VPWR 
+ VPWR
+ _4016_ sky130_fd_sc_hd__o21ai_1
X_8389_ _3605_ VGND VGND VPWR VPWR _4017_ sky130_fd_sc_hd__inv_2
X_8390_ _4017_ _3742_ VGND VGND VPWR VPWR 
+ _4018_
+ sky130_fd_sc_hd__or2_1
X_8391_ _4018_ VGND VGND VPWR VPWR _4019_ sky130_fd_sc_hd__clkinv_4
X_8392_ _3682_ VGND VGND VPWR VPWR _4020_ sky130_fd_sc_hd__inv_2
X_8393_ _3747_ VGND VGND VPWR VPWR _4021_ sky130_fd_sc_hd__inv_2
X_8394_ _3393_ _3383_ net142 _3390_ VGND VGND 
+ VPWR
+ VPWR _4022_ sky130_fd_sc_hd__or4_2
X_8395_ _3465_ _4022_ VGND VGND VPWR VPWR 
+ _4023_
+ sky130_fd_sc_hd__or2_1
X_8396_ _3800_ VGND VGND VPWR VPWR _4024_ sky130_fd_sc_hd__inv_2
X_8397_ _3513_ _3750_ VGND VGND VPWR VPWR 
+ _4025_
+ sky130_fd_sc_hd__nor2_1
X_8398_ _4024_ _4025_ _3751_ VGND VGND VPWR 
+ VPWR
+ _4026_ sky130_fd_sc_hd__o21ai_1
X_8399_ _3730_ _3746_ _4023_ _4026_ VGND VGND 
+ VPWR
+ VPWR _4027_ sky130_fd_sc_hd__o211a_1
X_8400_ _3437_ _3630_ _4021_ _4019_ _4027_ VGND 
+ VGND
+ VPWR VPWR _4028_ sky130_fd_sc_hd__o221a_1
X_8401_ _3628_ _4019_ VGND VGND VPWR VPWR 
+ _4029_
+ sky130_fd_sc_hd__or2_1
X_8402_ _3730_ _3630_ _3647_ _4028_ _4029_ VGND 
+ VGND
+ VPWR VPWR _4030_ sky130_fd_sc_hd__o2111a_1
X_8403_ _3651_ VGND VGND VPWR VPWR _4031_ sky130_fd_sc_hd__inv_2
X_8404_ _4031_ _3755_ VGND VGND VPWR VPWR 
+ _4032_
+ sky130_fd_sc_hd__or2_1
X_8405_ _4032_ VGND VGND VPWR VPWR _4033_ sky130_fd_sc_hd__inv_2
X_8406_ _3626_ _4019_ _4030_ _4033_ VGND VGND 
+ VPWR
+ VPWR _4034_ sky130_fd_sc_hd__o211a_1
X_8407_ _3654_ VGND VGND VPWR VPWR _4035_ sky130_fd_sc_hd__inv_2
X_8408_ _4035_ _3760_ VGND VGND VPWR VPWR 
+ _4036_
+ sky130_fd_sc_hd__nor2_1
X_8409_ _3623_ _4019_ _4034_ _4036_ VGND VGND 
+ VPWR
+ VPWR _4037_ sky130_fd_sc_hd__o211a_1
X_8410_ _3658_ VGND VGND VPWR VPWR _4038_ sky130_fd_sc_hd__inv_2
X_8411_ _4038_ _3767_ VGND VGND VPWR VPWR 
+ _4039_
+ sky130_fd_sc_hd__nor2_1
X_8412_ _3621_ _4019_ _4037_ _4039_ VGND VGND 
+ VPWR
+ VPWR _4040_ sky130_fd_sc_hd__o211a_1
X_8413_ _3662_ _3772_ VGND VGND VPWR VPWR 
+ _4041_
+ sky130_fd_sc_hd__or2_1
X_8414_ _4041_ VGND VGND VPWR VPWR _4042_ sky130_fd_sc_hd__inv_2
X_8415_ _3616_ _4019_ _4040_ _4042_ VGND VGND 
+ VPWR
+ VPWR _4043_ sky130_fd_sc_hd__o211a_1
X_8416_ _3668_ VGND VGND VPWR VPWR _4044_ sky130_fd_sc_hd__inv_2
X_8417_ _4044_ _3777_ VGND VGND VPWR VPWR 
+ _4045_
+ sky130_fd_sc_hd__or2_1
X_8418_ _4045_ VGND VGND VPWR VPWR _4046_ sky130_fd_sc_hd__inv_2
X_8419_ _3612_ _4019_ _4043_ _4046_ VGND VGND 
+ VPWR
+ VPWR _4047_ sky130_fd_sc_hd__o211a_1
X_8420_ _3674_ _3785_ VGND VGND VPWR VPWR 
+ _4048_
+ sky130_fd_sc_hd__or2_1
X_8421_ _4048_ VGND VGND VPWR VPWR _4049_ sky130_fd_sc_hd__inv_2
X_8422_ _3603_ _4019_ _4047_ _4049_ VGND VGND 
+ VPWR
+ VPWR _4050_ sky130_fd_sc_hd__o211a_1
X_8423_ _4020_ _3740_ _4050_ VGND VGND VPWR 
+ VPWR
+ _4051_ sky130_fd_sc_hd__or3b_1
X_8424_ _3681_ _4019_ _4051_ VGND VGND VPWR 
+ VPWR
+ _4052_ sky130_fd_sc_hd__o21bai_1
X_8425_ _3728_ _4016_ _4052_ VGND VGND VPWR 
+ VPWR
+ _4053_ sky130_fd_sc_hd__or3_1
X_8426_ _3458_ _3696_ VGND VGND VPWR VPWR 
+ _4054_
+ sky130_fd_sc_hd__or2_2
X_8427_ _4053_ _4054_ VGND VGND VPWR VPWR 
+ _4055_
+ sky130_fd_sc_hd__or2_1
X_8428_ _4015_ _4055_ VGND VGND VPWR VPWR 
+ _4056_
+ sky130_fd_sc_hd__or2_1
X_8429_ _3453_ _3585_ VGND VGND VPWR VPWR 
+ _4057_
+ sky130_fd_sc_hd__or2_1
X_8430_ _4056_ _4057_ VGND VGND VPWR VPWR 
+ _4058_
+ sky130_fd_sc_hd__or2_1
X_8431_ _3723_ _4058_ VGND VGND VPWR VPWR 
+ _4059_
+ sky130_fd_sc_hd__or2_1
X_8432_ _3434_ _3816_ _4059_ VGND VGND VPWR 
+ VPWR
+ _4060_ sky130_fd_sc_hd__or3_1
X_8433_ _3815_ _3718_ VGND VGND VPWR VPWR 
+ _4061_
+ sky130_fd_sc_hd__or2_1
X_8434_ _4060_ _4061_ VGND VGND VPWR VPWR 
+ _4062_
+ sky130_fd_sc_hd__nor2_1
X_8435_ _3813_ _4062_ VGND VGND VPWR VPWR 
+ _4063_
+ sky130_fd_sc_hd__or2_1
X_8436_ _4013_ _4063_ VGND VGND VPWR VPWR 
+ _4064_
+ sky130_fd_sc_hd__nand2_1
X_8437_ _3435_ _3582_ VGND VGND VPWR VPWR 
+ _4065_
+ sky130_fd_sc_hd__nor2_1
X_8438_ _3456_ _3481_ VGND VGND VPWR VPWR 
+ _4066_
+ sky130_fd_sc_hd__nor2_1
X_8439_ _3693_ _3689_ _3690_ _3691_ VGND VGND 
+ VPWR
+ VPWR _4067_ sky130_fd_sc_hd__a31o_1
X_8440_ _3495_ _3506_ _3613_ _3745_ VGND VGND 
+ VPWR
+ VPWR _4068_ sky130_fd_sc_hd__a2bb2o_1
X_8441_ _3522_ _3648_ VGND VGND VPWR VPWR 
+ _4069_
+ sky130_fd_sc_hd__nand2_1
X_8442_ _3519_ _3535_ _3433_ _3642_ VGND VGND 
+ VPWR
+ VPWR _4070_ sky130_fd_sc_hd__o22ai_1
X_8443_ _3532_ _3433_ _3527_ VGND VGND VPWR 
+ VPWR
+ _4071_ sky130_fd_sc_hd__o21ai_1
X_8444_ _4070_ _4071_ VGND VGND VPWR VPWR 
+ _4072_
+ sky130_fd_sc_hd__or2_1
X_8445_ _3452_ _3481_ _3584_ _3529_ _3426_ VGND 
+ VGND
+ VPWR VPWR _4073_ sky130_fd_sc_hd__a311o_1
X_8446_ _3495_ _3526_ _3639_ _4073_ _3643_ VGND 
+ VGND
+ VPWR VPWR _4074_ sky130_fd_sc_hd__o2111ai_2
X_8447_ _3465_ _3934_ VGND VGND VPWR VPWR 
+ _4075_
+ sky130_fd_sc_hd__or2_1
X_8448_ _3631_ _4072_ _4074_ _4075_ VGND VGND 
+ VPWR
+ VPWR _4076_ sky130_fd_sc_hd__or4b_1
X_8449_ _4069_ _4076_ VGND VGND VPWR VPWR 
+ _4077_
+ sky130_fd_sc_hd__or2_1
X_8450_ _3652_ VGND VGND VPWR VPWR _4078_ sky130_fd_sc_hd__inv_2
X_8451_ _3932_ _4078_ VGND VGND VPWR VPWR 
+ _4079_
+ sky130_fd_sc_hd__or2_1
X_8452_ _3504_ _3495_ _3446_ _3626_ VGND VGND 
+ VPWR
+ VPWR _4080_ sky130_fd_sc_hd__o22ai_1
X_8453_ _4068_ _4077_ _4079_ _4080_ VGND VGND 
+ VPWR
+ VPWR _4081_ sky130_fd_sc_hd__or4_1
X_8454_ _3542_ _3655_ VGND VGND VPWR VPWR 
+ _4082_
+ sky130_fd_sc_hd__nand2_1
X_8455_ _4081_ _4082_ VGND VGND VPWR VPWR 
+ _4083_
+ sky130_fd_sc_hd__or2_1
X_8456_ _3495_ _3499_ _3446_ _3623_ VGND VGND 
+ VPWR
+ VPWR _4084_ sky130_fd_sc_hd__o22ai_1
X_8457_ _3481_ _3501_ _3659_ VGND VGND VPWR 
+ VPWR
+ _4085_ sky130_fd_sc_hd__o21ai_2
X_8458_ _3495_ _3497_ _3446_ _3621_ VGND VGND 
+ VPWR
+ VPWR _4086_ sky130_fd_sc_hd__o22ai_1
X_8459_ _4083_ _4084_ _4085_ _4086_ VGND VGND 
+ VPWR
+ VPWR _4087_ sky130_fd_sc_hd__or4_1
X_8460_ _3664_ VGND VGND VPWR VPWR _4088_ sky130_fd_sc_hd__inv_2
X_8461_ _3949_ _4088_ VGND VGND VPWR VPWR 
+ _4089_
+ sky130_fd_sc_hd__or2_1
X_8462_ _3466_ _3492_ _3493_ _3613_ _3617_ VGND 
+ VGND
+ VPWR VPWR _4090_ sky130_fd_sc_hd__a32o_1
X_8463_ _3490_ _3670_ VGND VGND VPWR VPWR 
+ _4091_
+ sky130_fd_sc_hd__or2_1
X_8464_ _4087_ _4089_ _4090_ _4091_ VGND VGND 
+ VPWR
+ VPWR _4092_ sky130_fd_sc_hd__or4_1
X_8465_ _3476_ _3483_ _3446_ _3612_ VGND VGND 
+ VPWR
+ VPWR _4093_ sky130_fd_sc_hd__o22ai_1
X_8466_ _4092_ _4093_ VGND VGND VPWR VPWR 
+ _4094_
+ sky130_fd_sc_hd__or2_1
X_8467_ _3676_ VGND VGND VPWR VPWR _4095_ sky130_fd_sc_hd__inv_2
X_8468_ _3954_ _4095_ VGND VGND VPWR VPWR 
+ _4096_
+ sky130_fd_sc_hd__or2_1
X_8469_ _3473_ _3476_ _3446_ _3603_ VGND VGND 
+ VPWR
+ VPWR _4097_ sky130_fd_sc_hd__o22ai_1
X_8470_ _4094_ _4096_ _4097_ VGND VGND VPWR 
+ VPWR
+ _4098_ sky130_fd_sc_hd__or3_1
X_8471_ _3421_ VGND VGND VPWR VPWR _4099_ sky130_fd_sc_hd__clkinv_2
X_8472_ _3530_ VGND VGND VPWR VPWR _4100_ sky130_fd_sc_hd__clkinv_2
X_8473_ _4099_ _4100_ _3688_ _3684_ VGND VGND 
+ VPWR
+ VPWR _4101_ sky130_fd_sc_hd__a31o_1
X_8474_ _4098_ _4101_ VGND VGND VPWR VPWR 
+ _4102_
+ sky130_fd_sc_hd__or2_1
X_8475_ _3694_ _4067_ _4102_ VGND VGND VPWR 
+ VPWR
+ _4103_ sky130_fd_sc_hd__or3_1
X_8476_ _3458_ _3833_ VGND VGND VPWR VPWR 
+ _4104_
+ sky130_fd_sc_hd__or2_2
X_8477_ _4103_ _4104_ VGND VGND VPWR VPWR 
+ _4105_
+ sky130_fd_sc_hd__or2_1
X_8478_ _4066_ _4105_ VGND VGND VPWR VPWR 
+ _4106_
+ sky130_fd_sc_hd__or2_1
X_8479_ _4065_ _4106_ VGND VGND VPWR VPWR 
+ _4107_
+ sky130_fd_sc_hd__or2_1
X_8480_ _3472_ _3582_ _3481_ _3582_ VGND VGND 
+ VPWR
+ VPWR _4108_ sky130_fd_sc_hd__o22ai_4
X_8481_ _4107_ _4108_ VGND VGND VPWR VPWR 
+ _4109_
+ sky130_fd_sc_hd__or2_1
X_8482_ _3434_ _3817_ VGND VGND VPWR VPWR 
+ _4110_
+ sky130_fd_sc_hd__or2_1
X_8483_ _4109_ _4110_ VGND VGND VPWR VPWR 
+ _4111_
+ sky130_fd_sc_hd__or2_1
X_8484_ _3428_ _3605_ _3715_ VGND VGND VPWR 
+ VPWR
+ _4112_ sky130_fd_sc_hd__o21ai_1
X_8485_ _4111_ _4112_ VGND VGND VPWR VPWR 
+ _4113_
+ sky130_fd_sc_hd__or2_1
X_8486_ _3575_ _4113_ VGND VGND VPWR VPWR 
+ _4114_
+ sky130_fd_sc_hd__or2b_1
X_8487_ _4064_ _4114_ VGND VGND VPWR VPWR 
+ _4115_
+ sky130_fd_sc_hd__or2b_1
X_8488_ _4115_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
X_8489_ _3724_ _3701_ _3453_ VGND VGND VPWR 
+ VPWR
+ _4116_ sky130_fd_sc_hd__or3_1
X_8490_ _3502_ _3876_ _3945_ VGND VGND VPWR 
+ VPWR
+ _4117_ sky130_fd_sc_hd__or3_1
X_8491_ _3493_ _3931_ _3491_ _3892_ VGND VGND 
+ VPWR
+ VPWR _4118_ sky130_fd_sc_hd__a211o_1
X_8492_ _3549_ VGND VGND VPWR VPWR _4119_ sky130_fd_sc_hd__inv_2
X_8493_ _4119_ _3884_ _3948_ VGND VGND VPWR 
+ VPWR
+ _4120_ sky130_fd_sc_hd__or3_1
X_8494_ _3472_ _3476_ _3385_ _3465_ _3526_ VGND 
+ VGND
+ VPWR VPWR _4121_ sky130_fd_sc_hd__a311oi_2
X_8495_ _3444_ _3535_ _3396_ _3516_ VGND VGND 
+ VPWR
+ VPWR _4122_ sky130_fd_sc_hd__o22a_1
X_8496_ _3465_ _4122_ VGND VGND VPWR VPWR 
+ _4123_
+ sky130_fd_sc_hd__nor2_2
X_8497_ _3937_ _4023_ VGND VGND VPWR VPWR 
+ _4124_
+ sky130_fd_sc_hd__or2b_1
X_8498_ _3535_ _3930_ VGND VGND VPWR VPWR 
+ _4125_
+ sky130_fd_sc_hd__nor2_1
X_8499_ _3855_ _3856_ VGND VGND VPWR VPWR 
+ _4126_
+ sky130_fd_sc_hd__or2_1
X_8500_ _4125_ _4126_ _3969_ _3523_ VGND VGND 
+ VPWR
+ VPWR _4127_ sky130_fd_sc_hd__or4b_1
X_8501_ _4121_ _4123_ _4124_ _4127_ VGND VGND 
+ VPWR
+ VPWR _4128_ sky130_fd_sc_hd__or4_2
X_8502_ _3506_ _3930_ _3508_ _3862_ VGND VGND 
+ VPWR
+ VPWR _4129_ sky130_fd_sc_hd__o211a_1
X_8503_ _3444_ _3505_ _3504_ _3930_ _3541_ VGND 
+ VGND
+ VPWR VPWR _4130_ sky130_fd_sc_hd__o221a_1
X_8504_ _4128_ _4129_ _4130_ VGND VGND VPWR 
+ VPWR
+ _4131_ sky130_fd_sc_hd__and3b_1
X_8505_ _4117_ _4118_ _4120_ _4131_ VGND VGND 
+ VPWR
+ VPWR _4132_ sky130_fd_sc_hd__or4b_4
X_8506_ _3485_ _3900_ _3953_ VGND VGND VPWR 
+ VPWR
+ _4133_ sky130_fd_sc_hd__or3_2
X_8507_ _3468_ _3511_ _3473_ _3928_ _3474_ VGND 
+ VGND
+ VPWR VPWR _4134_ sky130_fd_sc_hd__o221ai_2
X_8508_ _3389_ _3462_ _3393_ _3397_ _3959_ VGND 
+ VGND
+ VPWR VPWR _4135_ sky130_fd_sc_hd__a41o_1
X_8509_ _4132_ _4133_ _4134_ _4135_ VGND VGND 
+ VPWR
+ VPWR _4136_ sky130_fd_sc_hd__or4_1
X_8510_ _3395_ _3450_ _3388_ VGND VGND VPWR 
+ VPWR
+ _4137_ sky130_fd_sc_hd__nor3_1
X_8511_ _3389_ _3635_ _3439_ _3926_ VGND VGND 
+ VPWR
+ VPWR _4138_ sky130_fd_sc_hd__a211o_1
X_8512_ _4116_ _4136_ _4137_ _4138_ VGND VGND 
+ VPWR
+ VPWR _4139_ sky130_fd_sc_hd__or4_1
X_8513_ _4139_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
X_8514_ _3815_ _3575_ _4112_ VGND VGND VPWR 
+ VPWR
+ _4140_ sky130_fd_sc_hd__or3_1
X_8515_ _3456_ _3472_ VGND VGND VPWR VPWR 
+ _4141_
+ sky130_fd_sc_hd__nor2_1
X_8516_ _3529_ _3425_ VGND VGND VPWR VPWR 
+ _4142_
+ sky130_fd_sc_hd__nor2_4
X_8517_ _3531_ VGND VGND VPWR VPWR _4143_ sky130_fd_sc_hd__inv_2
X_8518_ _3693_ _4017_ VGND VGND VPWR VPWR 
+ _4144_
+ sky130_fd_sc_hd__or2_4
X_8519_ _4142_ _4143_ _4144_ _4079_ VGND VGND 
+ VPWR
+ VPWR _4145_ sky130_fd_sc_hd__a31o_1
X_8520_ _4100_ _4143_ _4144_ _4071_ VGND VGND 
+ VPWR
+ VPWR _4146_ sky130_fd_sc_hd__a31o_1
X_8521_ _3437_ _3481_ VGND VGND VPWR VPWR 
+ _4147_
+ sky130_fd_sc_hd__nand2_1
X_8522_ _3636_ _3689_ _4147_ _3640_ VGND VGND 
+ VPWR
+ VPWR _4148_ sky130_fd_sc_hd__a31o_1
X_8523_ _3641_ VGND VGND VPWR VPWR _4149_ sky130_fd_sc_hd__inv_2
X_8524_ _4149_ _4143_ _4144_ _4070_ VGND VGND 
+ VPWR
+ VPWR _4150_ sky130_fd_sc_hd__a31o_1
X_8525_ net158 _3424_ _3529_ VGND VGND VPWR 
+ VPWR
+ _4151_ sky130_fd_sc_hd__nor3_4
X_8526_ _4151_ _4143_ _4144_ _4069_ VGND VGND 
+ VPWR
+ VPWR _4152_ sky130_fd_sc_hd__a31o_1
X_8527_ _4146_ _4148_ _4150_ _4152_ VGND VGND 
+ VPWR
+ VPWR _4153_ sky130_fd_sc_hd__or4_1
X_8528_ net160 _3419_ VGND VGND VPWR VPWR 
+ _4154_
+ sky130_fd_sc_hd__nor2_4
X_8529_ _4149_ _4154_ _4144_ _4082_ VGND VGND 
+ VPWR
+ VPWR _4155_ sky130_fd_sc_hd__a31o_1
X_8530_ _4100_ _4154_ _4144_ _4085_ VGND VGND 
+ VPWR
+ VPWR _4156_ sky130_fd_sc_hd__a31o_1
X_8531_ _4145_ _4153_ _4155_ _4156_ VGND VGND 
+ VPWR
+ VPWR _4157_ sky130_fd_sc_hd__or4_1
X_8532_ _4154_ _4151_ _4144_ _4089_ VGND VGND 
+ VPWR
+ VPWR _4158_ sky130_fd_sc_hd__a31o_1
X_8533_ _4142_ _4154_ _4144_ _4091_ VGND VGND 
+ VPWR
+ VPWR _4159_ sky130_fd_sc_hd__a31o_1
X_8534_ _4099_ _4149_ _4144_ _4096_ VGND VGND 
+ VPWR
+ VPWR _4160_ sky130_fd_sc_hd__a31o_1
X_8535_ _4157_ _4158_ _4159_ _4160_ VGND VGND 
+ VPWR
+ VPWR _4161_ sky130_fd_sc_hd__or4_2
X_8536_ _3686_ VGND VGND VPWR VPWR _4162_ sky130_fd_sc_hd__inv_2
X_8537_ _3391_ _3492_ _3690_ _4162_ _4101_ VGND 
+ VGND
+ VPWR VPWR _4163_ sky130_fd_sc_hd__a311o_1
X_8538_ _3404_ _3424_ _3421_ _3714_ VGND VGND 
+ VPWR
+ VPWR _4164_ sky130_fd_sc_hd__or4_1
X_8539_ _3696_ _4104_ _4164_ VGND VGND VPWR 
+ VPWR
+ _4165_ sky130_fd_sc_hd__or3b_2
X_8540_ _3702_ _4065_ VGND VGND VPWR VPWR 
+ _4166_
+ sky130_fd_sc_hd__or2_1
X_8541_ _4161_ _4163_ _4165_ _4166_ VGND VGND 
+ VPWR
+ VPWR _4167_ sky130_fd_sc_hd__nor4_1
X_8542_ _4141_ _4110_ _3967_ _4167_ VGND VGND 
+ VPWR
+ VPWR _4168_ sky130_fd_sc_hd__or4b_1
X_8543_ _4168_ VGND VGND VPWR VPWR _4169_ sky130_fd_sc_hd__inv_2
X_8544_ _3613_ _3741_ _4018_ VGND VGND VPWR 
+ VPWR
+ _4170_ sky130_fd_sc_hd__or3_2
X_8545_ _4170_ VGND VGND VPWR VPWR _4171_ sky130_fd_sc_hd__clkinv_4
X_8546_ _3749_ _3635_ VGND VGND VPWR VPWR 
+ _4172_
+ sky130_fd_sc_hd__nor2_1
X_8547_ _3600_ _4172_ _4026_ VGND VGND VPWR 
+ VPWR
+ _4173_ sky130_fd_sc_hd__o21a_1
X_8548_ _4021_ _4171_ _3628_ _4171_ _4173_ VGND 
+ VGND
+ VPWR VPWR _4174_ sky130_fd_sc_hd__o221a_1
X_8549_ _3626_ _4171_ _3623_ _4171_ _4174_ VGND 
+ VGND
+ VPWR VPWR _4175_ sky130_fd_sc_hd__o221ai_1
X_8550_ _3621_ _4171_ VGND VGND VPWR VPWR 
+ _4176_
+ sky130_fd_sc_hd__nor2_1
X_8551_ _3616_ _4171_ VGND VGND VPWR VPWR 
+ _4177_
+ sky130_fd_sc_hd__nor2_1
X_8552_ _3612_ _4171_ VGND VGND VPWR VPWR 
+ _4178_
+ sky130_fd_sc_hd__nor2_1
X_8553_ _4175_ _4176_ _4177_ _4178_ VGND VGND 
+ VPWR
+ VPWR _4179_ sky130_fd_sc_hd__or4_2
X_8554_ _3603_ _4171_ VGND VGND VPWR VPWR 
+ _4180_
+ sky130_fd_sc_hd__nor2_1
X_8555_ _3438_ _3750_ _3681_ _4019_ _3798_ VGND 
+ VGND
+ VPWR VPWR _4181_ sky130_fd_sc_hd__o221ai_1
X_8556_ _4054_ VGND VGND VPWR VPWR _4182_ sky130_fd_sc_hd__inv_2
X_8557_ _3720_ _3595_ _3605_ _3459_ _4182_ VGND 
+ VGND
+ VPWR VPWR _4183_ sky130_fd_sc_hd__o311a_1
X_8558_ _4183_ VGND VGND VPWR VPWR _4184_ sky130_fd_sc_hd__inv_2
X_8559_ _4179_ _4180_ _4181_ _4184_ VGND VGND 
+ VPWR
+ VPWR _4185_ sky130_fd_sc_hd__or4_1
X_8560_ _3725_ _4057_ VGND VGND VPWR VPWR 
+ _4186_
+ sky130_fd_sc_hd__or2_2
X_8561_ _3433_ _4014_ VGND VGND VPWR VPWR 
+ _4187_
+ sky130_fd_sc_hd__nor2_1
X_8562_ _3434_ _3816_ _3926_ VGND VGND VPWR 
+ VPWR
+ _4188_ sky130_fd_sc_hd__or3_1
X_8563_ _4185_ _4186_ _4187_ _4188_ VGND VGND 
+ VPWR
+ VPWR _4189_ sky130_fd_sc_hd__or4_1
X_8564_ _3392_ _3813_ _4061_ _4189_ VGND VGND 
+ VPWR
+ VPWR _4190_ sky130_fd_sc_hd__or4b_1
X_8565_ _4005_ _3710_ VGND VGND VPWR VPWR 
+ _4191_
+ sky130_fd_sc_hd__nor2_1
X_8566_ _3512_ _3635_ VGND VGND VPWR VPWR 
+ _4192_
+ sky130_fd_sc_hd__nor2_1
X_8567_ _3738_ _4192_ _3972_ VGND VGND VPWR 
+ VPWR
+ _4193_ sky130_fd_sc_hd__o21ai_2
X_8568_ _3730_ _3978_ _3845_ VGND VGND VPWR 
+ VPWR
+ _4194_ sky130_fd_sc_hd__o21a_1
X_8569_ _3738_ _4194_ _3851_ _3979_ VGND VGND 
+ VPWR
+ VPWR _4195_ sky130_fd_sc_hd__o211ai_4
X_8570_ _3730_ _3630_ _3526_ _3840_ _3977_ VGND 
+ VGND
+ VPWR VPWR _4196_ sky130_fd_sc_hd__o221ai_4
X_8571_ _3755_ _3855_ _3982_ VGND VGND VPWR 
+ VPWR
+ _4197_ sky130_fd_sc_hd__or3_1
X_8572_ _4193_ _4195_ _4196_ _4197_ VGND VGND 
+ VPWR
+ VPWR _4198_ sky130_fd_sc_hd__or4_1
X_8573_ _3760_ _3860_ _3985_ VGND VGND VPWR 
+ VPWR
+ _4199_ sky130_fd_sc_hd__or3_1
X_8574_ _3767_ _3868_ _3987_ VGND VGND VPWR 
+ VPWR
+ _4200_ sky130_fd_sc_hd__or3_1
X_8575_ _3772_ _3874_ _3990_ VGND VGND VPWR 
+ VPWR
+ _4201_ sky130_fd_sc_hd__or3_1
X_8576_ _4198_ _4199_ _4200_ _4201_ VGND VGND 
+ VPWR
+ VPWR _4202_ sky130_fd_sc_hd__or4_1
X_8577_ _3777_ _3882_ _3993_ VGND VGND VPWR 
+ VPWR
+ _4203_ sky130_fd_sc_hd__or3_1
X_8578_ _3785_ _3890_ _3995_ VGND VGND VPWR 
+ VPWR
+ _4204_ sky130_fd_sc_hd__or3_1
X_8579_ _3740_ _3898_ _3998_ VGND VGND VPWR 
+ VPWR
+ _4205_ sky130_fd_sc_hd__or3_2
X_8580_ _4202_ _4203_ _4204_ _4205_ VGND VGND 
+ VPWR
+ VPWR _4206_ sky130_fd_sc_hd__or4_4
X_8581_ _3634_ _3848_ _3906_ VGND VGND VPWR 
+ VPWR
+ _4207_ sky130_fd_sc_hd__o21ai_1
X_8582_ _4001_ _4207_ VGND VGND VPWR VPWR 
+ _4208_
+ sky130_fd_sc_hd__or2_1
X_8583_ _3404_ _3821_ _3827_ VGND VGND VPWR 
+ VPWR
+ _4209_ sky130_fd_sc_hd__nor3_1
X_8584_ _3831_ _3741_ _4209_ _3912_ _4004_ VGND 
+ VGND
+ VPWR VPWR _4210_ sky130_fd_sc_hd__a311o_1
X_8585_ _4007_ _3585_ VGND VGND VPWR VPWR 
+ _4211_
+ sky130_fd_sc_hd__or2_1
X_8586_ _4206_ _4208_ _4210_ _4211_ VGND VGND 
+ VPWR
+ VPWR _4212_ sky130_fd_sc_hd__or4_1
X_8587_ _3439_ _3818_ VGND VGND VPWR VPWR 
+ _4213_
+ sky130_fd_sc_hd__or2_1
X_8588_ _4191_ _4212_ _3967_ _4213_ VGND VGND 
+ VPWR
+ VPWR _4214_ sky130_fd_sc_hd__or4_1
X_8589_ _3817_ _3923_ _4011_ _4214_ VGND VGND 
+ VPWR
+ VPWR _4215_ sky130_fd_sc_hd__or4b_2
X_8590_ _4140_ _4169_ _4190_ _4215_ VGND VGND 
+ VPWR
+ VPWR _0183_ sky130_fd_sc_hd__o211ai_1
X_8591_ _3395_ _3535_ _3509_ _3513_ VGND VGND 
+ VPWR
+ VPWR _4216_ sky130_fd_sc_hd__o211ai_1
X_8592_ _3940_ VGND VGND VPWR VPWR _4217_ sky130_fd_sc_hd__inv_2
X_8593_ _3466_ _4216_ _4217_ _4124_ VGND VGND 
+ VPWR
+ VPWR _4218_ sky130_fd_sc_hd__a211o_1
X_8594_ _4121_ _3969_ _3527_ VGND VGND VPWR 
+ VPWR
+ _4219_ sky130_fd_sc_hd__or3b_1
X_8595_ _4219_ _3835_ _3838_ _3533_ VGND VGND 
+ VPWR
+ VPWR _4220_ sky130_fd_sc_hd__or4b_1
X_8596_ _3478_ _3505_ _3865_ _3933_ _4129_ VGND 
+ VGND
+ VPWR VPWR _4221_ sky130_fd_sc_hd__o2111ai_4
X_8597_ _3547_ _3880_ _3946_ _4117_ VGND VGND 
+ VPWR
+ VPWR _4222_ sky130_fd_sc_hd__or4_4
X_8598_ _4218_ _4220_ _4221_ _4222_ VGND VGND 
+ VPWR
+ VPWR _4223_ sky130_fd_sc_hd__or4_2
X_8599_ _3486_ _3896_ _3952_ _4118_ VGND VGND 
+ VPWR
+ VPWR _4224_ sky130_fd_sc_hd__or4_4
X_8600_ _3927_ _4134_ VGND VGND VPWR VPWR 
+ _4225_
+ sky130_fd_sc_hd__or2_1
X_8601_ _4223_ _4224_ _4225_ _4054_ VGND VGND 
+ VPWR
+ VPWR _4226_ sky130_fd_sc_hd__or4_1
X_8602_ _3442_ _3444_ _3388_ _3511_ _3963_ VGND 
+ VGND
+ VPWR VPWR _4227_ sky130_fd_sc_hd__o221ai_1
X_8603_ _4116_ _4226_ _4137_ _4227_ VGND VGND 
+ VPWR
+ VPWR _4228_ sky130_fd_sc_hd__or4_1
X_8604_ _4228_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_8605_ _4110_ _4140_ VGND VGND VPWR VPWR 
+ _4229_
+ sky130_fd_sc_hd__or2_1
X_8606_ _3707_ _3818_ VGND VGND VPWR VPWR 
+ _4230_
+ sky130_fd_sc_hd__or2_1
X_8607_ _4145_ _4035_ _4080_ _3541_ VGND VGND 
+ VPWR
+ VPWR _4231_ sky130_fd_sc_hd__or4b_2
X_8608_ _3465_ _3472_ _3521_ _3647_ _4075_ VGND 
+ VGND
+ VPWR VPWR _4232_ sky130_fd_sc_hd__o311a_1
X_8609_ _4232_ VGND VGND VPWR VPWR _4233_ sky130_fd_sc_hd__inv_2
X_8610_ _3396_ _3516_ _3511_ VGND VGND VPWR 
+ VPWR
+ _4234_ sky130_fd_sc_hd__o21ai_1
X_8611_ _3636_ _4234_ _3637_ _4148_ VGND VGND 
+ VPWR
+ VPWR _4235_ sky130_fd_sc_hd__a211o_1
X_8612_ _3631_ _4146_ VGND VGND VPWR VPWR 
+ _4236_
+ sky130_fd_sc_hd__or2_1
X_8613_ _4233_ _4235_ _4236_ VGND VGND VPWR 
+ VPWR
+ _4237_ sky130_fd_sc_hd__or3_1
X_8614_ _4119_ _3662_ _4086_ _4156_ VGND VGND 
+ VPWR
+ VPWR _4238_ sky130_fd_sc_hd__or4_1
X_8615_ _3485_ _3674_ _4093_ _4159_ VGND VGND 
+ VPWR
+ VPWR _4239_ sky130_fd_sc_hd__or4_1
X_8616_ _4231_ _4237_ _4238_ _4239_ VGND VGND 
+ VPWR
+ VPWR _4240_ sky130_fd_sc_hd__or4_2
X_8617_ _4067_ _4163_ VGND VGND VPWR VPWR 
+ _4241_
+ sky130_fd_sc_hd__or2_1
X_8618_ _3456_ _3476_ _3437_ _3456_ VGND VGND 
+ VPWR
+ VPWR _4242_ sky130_fd_sc_hd__o22ai_2
X_8619_ _4240_ _4241_ _4242_ _4166_ VGND VGND 
+ VPWR
+ VPWR _4243_ sky130_fd_sc_hd__or4_1
X_8620_ _4108_ _4230_ _4141_ _4243_ VGND VGND 
+ VPWR
+ VPWR _4244_ sky130_fd_sc_hd__nor4_1
X_8621_ _4186_ VGND VGND VPWR VPWR _4245_ sky130_fd_sc_hd__inv_2
X_8622_ _3595_ _3624_ _3433_ _3513_ _4022_ VGND 
+ VGND
+ VPWR VPWR _4246_ sky130_fd_sc_hd__o311a_1
X_8623_ _3600_ _4246_ _4173_ VGND VGND VPWR 
+ VPWR
+ _4247_ sky130_fd_sc_hd__o21ai_2
X_8624_ _3435_ _3433_ VGND VGND VPWR VPWR 
+ _4248_
+ sky130_fd_sc_hd__and2_1
X_8625_ _3731_ _4170_ VGND VGND VPWR VPWR 
+ _4249_
+ sky130_fd_sc_hd__nor2_1
X_8626_ _3628_ _4248_ _3630_ _4249_ VGND VGND 
+ VPWR
+ VPWR _4250_ sky130_fd_sc_hd__o22ai_2
X_8627_ _4088_ _3773_ _4041_ _4176_ VGND VGND 
+ VPWR
+ VPWR _4251_ sky130_fd_sc_hd__or4_2
X_8628_ _3626_ _4171_ _3655_ _3762_ _4036_ VGND 
+ VGND
+ VPWR VPWR _4252_ sky130_fd_sc_hd__o2111a_1
X_8629_ _4247_ _4250_ _4251_ _4252_ VGND VGND 
+ VPWR
+ VPWR _4253_ sky130_fd_sc_hd__or4b_2
X_8630_ _4095_ _3787_ _4048_ _4178_ VGND VGND 
+ VPWR
+ VPWR _4254_ sky130_fd_sc_hd__or4_2
X_8631_ _4016_ _4181_ VGND VGND VPWR VPWR 
+ _4255_
+ sky130_fd_sc_hd__or2_1
X_8632_ _3435_ _4014_ VGND VGND VPWR VPWR 
+ _4256_
+ sky130_fd_sc_hd__nor2_1
X_8633_ _4253_ _4254_ _4255_ _4256_ VGND VGND 
+ VPWR
+ VPWR _4257_ sky130_fd_sc_hd__nor4_1
X_8634_ _3613_ _3722_ _3439_ _3723_ VGND VGND 
+ VPWR
+ VPWR _4258_ sky130_fd_sc_hd__a211o_1
X_8635_ _4187_ _4258_ VGND VGND VPWR VPWR 
+ _4259_
+ sky130_fd_sc_hd__nor2_1
X_8636_ _3392_ _3813_ _4061_ _4188_ VGND VGND 
+ VPWR
+ VPWR _4260_ sky130_fd_sc_hd__or4_2
X_8637_ _4245_ _4257_ _4259_ _4260_ VGND VGND 
+ VPWR
+ VPWR _4261_ sky130_fd_sc_hd__a31o_1
X_8638_ _4211_ VGND VGND VPWR VPWR _4262_ sky130_fd_sc_hd__inv_2
X_8639_ _3745_ _3742_ _3838_ _3970_ _4196_ VGND 
+ VGND
+ VPWR VPWR _4263_ sky130_fd_sc_hd__a2111o_1
X_8640_ _3738_ _3710_ _3978_ VGND VGND VPWR 
+ VPWR
+ _4264_ sky130_fd_sc_hd__nor3_1
X_8641_ _4217_ _4193_ _4264_ _3971_ VGND VGND 
+ VPWR
+ VPWR _4265_ sky130_fd_sc_hd__or4b_2
X_8642_ _3764_ _3864_ _3986_ _4199_ VGND VGND 
+ VPWR
+ VPWR _4266_ sky130_fd_sc_hd__or4_2
X_8643_ _3617_ _3742_ _3877_ _3991_ _4201_ VGND 
+ VGND
+ VPWR VPWR _4267_ sky130_fd_sc_hd__a2111o_2
X_8644_ _4263_ _4265_ _4266_ _4267_ VGND VGND 
+ VPWR
+ VPWR _4268_ sky130_fd_sc_hd__or4_4
X_8645_ _3789_ _3894_ _3997_ _4204_ VGND VGND 
+ VPWR
+ VPWR _4269_ sky130_fd_sc_hd__or4_4
X_8646_ _4002_ _4208_ VGND VGND VPWR VPWR 
+ _4270_
+ sky130_fd_sc_hd__or2_1
X_8647_ _4268_ _4269_ _4270_ _4104_ VGND VGND 
+ VPWR
+ VPWR _4271_ sky130_fd_sc_hd__nor4_1
X_8648_ _3635_ _3844_ _3831_ VGND VGND VPWR 
+ VPWR
+ _4272_ sky130_fd_sc_hd__o21a_1
X_8649_ _3968_ _4272_ _4191_ VGND VGND VPWR 
+ VPWR
+ _4273_ sky130_fd_sc_hd__nor3_1
X_8650_ _3816_ _3817_ _3923_ VGND VGND VPWR 
+ VPWR
+ _4274_ sky130_fd_sc_hd__or3_1
X_8651_ _3429_ _4011_ VGND VGND VPWR VPWR 
+ _4275_
+ sky130_fd_sc_hd__or2_1
X_8652_ _4213_ _4274_ _4275_ VGND VGND VPWR 
+ VPWR
+ _4276_ sky130_fd_sc_hd__or3_1
X_8653_ _4262_ _4271_ _4273_ _4276_ VGND VGND 
+ VPWR
+ VPWR _4277_ sky130_fd_sc_hd__a31o_1
X_8654_ _3967_ _4229_ _4244_ _4261_ _4277_ VGND 
+ VGND
+ VPWR VPWR _4278_ sky130_fd_sc_hd__o311a_1
X_8655_ _4278_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__inv_2
X_8656_ _3466_ _3493_ _3693_ _3888_ VGND VGND 
+ VPWR
+ VPWR _4279_ sky130_fd_sc_hd__a31o_1
X_8657_ _3950_ _4279_ _4120_ _4222_ VGND VGND 
+ VPWR
+ VPWR _4280_ sky130_fd_sc_hd__or4_2
X_8658_ _3858_ _3859_ VGND VGND VPWR VPWR 
+ _4281_
+ sky130_fd_sc_hd__or2_1
X_8659_ _4126_ _4281_ _4220_ _3524_ VGND VGND 
+ VPWR
+ VPWR _4282_ sky130_fd_sc_hd__or4b_1
X_8660_ _3385_ _3450_ _3388_ VGND VGND VPWR 
+ VPWR
+ _4283_ sky130_fd_sc_hd__or3_1
X_8661_ _3388_ _3444_ _3450_ _4283_ _4182_ VGND 
+ VGND
+ VPWR VPWR _4284_ sky130_fd_sc_hd__o311a_1
X_8662_ _3467_ _4135_ _4225_ _4284_ VGND VGND 
+ VPWR
+ VPWR _4285_ sky130_fd_sc_hd__or4b_2
X_8663_ _4280_ _4282_ _4285_ _3832_ VGND VGND 
+ VPWR
+ VPWR _4286_ sky130_fd_sc_hd__or4_1
X_8664_ _4286_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
X_8665_ _4068_ _4031_ _3508_ VGND VGND VPWR 
+ VPWR
+ _4287_ sky130_fd_sc_hd__or3b_1
X_8666_ _4152_ _4287_ _4233_ _4236_ VGND VGND 
+ VPWR
+ VPWR _4288_ sky130_fd_sc_hd__or4_2
X_8667_ _3491_ _4044_ VGND VGND VPWR VPWR 
+ _4289_
+ sky130_fd_sc_hd__or2_1
X_8668_ _4090_ _4289_ _4158_ _4238_ VGND VGND 
+ VPWR
+ VPWR _4290_ sky130_fd_sc_hd__or4_4
X_8669_ _3701_ _4066_ _4242_ VGND VGND VPWR 
+ VPWR
+ _4291_ sky130_fd_sc_hd__or3_1
X_8670_ _3694_ _4165_ _4291_ _4241_ VGND VGND 
+ VPWR
+ VPWR _4292_ sky130_fd_sc_hd__or4_1
X_8671_ _4288_ _4290_ _4292_ _3453_ VGND VGND 
+ VPWR
+ VPWR _4293_ sky130_fd_sc_hd__nor4_2
X_8672_ _4141_ _3707_ _3816_ VGND VGND VPWR 
+ VPWR
+ _4294_ sky130_fd_sc_hd__or3_1
X_8673_ _3926_ _4108_ _4294_ _4229_ VGND VGND 
+ VPWR
+ VPWR _4295_ sky130_fd_sc_hd__or4_2
X_8674_ _3781_ _3886_ VGND VGND VPWR VPWR 
+ _4296_
+ sky130_fd_sc_hd__or2_1
X_8675_ _3994_ _4296_ _4203_ _4267_ VGND VGND 
+ VPWR
+ VPWR _4297_ sky130_fd_sc_hd__or4_4
X_8676_ _3758_ _3858_ VGND VGND VPWR VPWR 
+ _4298_
+ sky130_fd_sc_hd__or2_1
X_8677_ _3983_ _4298_ _4197_ _4263_ VGND VGND 
+ VPWR
+ VPWR _4299_ sky130_fd_sc_hd__or4_4
X_8678_ _3834_ _4210_ _4270_ VGND VGND VPWR 
+ VPWR
+ _4300_ sky130_fd_sc_hd__or3_2
X_8679_ _3832_ _4006_ _4104_ _4300_ VGND VGND 
+ VPWR
+ VPWR _4301_ sky130_fd_sc_hd__or4_4
X_8680_ _4297_ _4299_ _4301_ _3724_ VGND VGND 
+ VPWR
+ VPWR _4302_ sky130_fd_sc_hd__nor4_2
X_8681_ _4213_ _4272_ _4275_ VGND VGND VPWR 
+ VPWR
+ _4303_ sky130_fd_sc_hd__or3_1
X_8682_ _4191_ _3968_ _4274_ _4303_ VGND VGND 
+ VPWR
+ VPWR _4304_ sky130_fd_sc_hd__or4_4
X_8683_ _4078_ _3756_ VGND VGND VPWR VPWR 
+ _4305_
+ sky130_fd_sc_hd__or2_1
X_8684_ _3745_ _4170_ _4032_ _4305_ _4250_ VGND 
+ VGND
+ VPWR VPWR _4306_ sky130_fd_sc_hd__a2111o_2
X_8685_ _3670_ _3779_ VGND VGND VPWR VPWR 
+ _4307_
+ sky130_fd_sc_hd__or2_1
X_8686_ _4045_ _4307_ _4177_ _4251_ VGND VGND 
+ VPWR
+ VPWR _4308_ sky130_fd_sc_hd__or4_2
X_8687_ _3724_ _4015_ _4256_ VGND VGND VPWR 
+ VPWR
+ _4309_ sky130_fd_sc_hd__or3_1
X_8688_ _3728_ _4184_ _4255_ VGND VGND VPWR 
+ VPWR
+ _4310_ sky130_fd_sc_hd__or3_1
X_8689_ _4306_ _4308_ _4309_ _4310_ VGND VGND 
+ VPWR
+ VPWR _4311_ sky130_fd_sc_hd__or4_1
X_8690_ _4260_ VGND VGND VPWR VPWR _4312_ sky130_fd_sc_hd__inv_2
X_8691_ _3701_ _4311_ _4259_ _4312_ VGND VGND 
+ VPWR
+ VPWR _4313_ sky130_fd_sc_hd__o211ai_2
X_8692_ _4293_ _4295_ _4302_ _4304_ _4313_ VGND 
+ VGND
+ VPWR VPWR _0187_ sky130_fd_sc_hd__o221ai_4
X_8693_ _4133_ _3904_ _3955_ _3479_ VGND VGND 
+ VPWR
+ VPWR _4314_ sky130_fd_sc_hd__or4b_1
X_8694_ _3465_ _3846_ _3841_ _3536_ VGND VGND 
+ VPWR
+ VPWR _4315_ sky130_fd_sc_hd__o211ai_1
X_8695_ _4125_ _4315_ _4123_ _4218_ VGND VGND 
+ VPWR
+ VPWR _4316_ sky130_fd_sc_hd__or4_1
X_8696_ _4224_ _4314_ _4280_ _4316_ VGND VGND 
+ VPWR
+ VPWR _4317_ sky130_fd_sc_hd__or4_1
X_8697_ _4317_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
X_8698_ _4097_ _4020_ _3474_ VGND VGND VPWR 
+ VPWR
+ _4318_ sky130_fd_sc_hd__or3b_1
X_8699_ _4160_ _4318_ _4239_ _4290_ VGND VGND 
+ VPWR
+ VPWR _4319_ sky130_fd_sc_hd__or4_1
X_8700_ _3472_ _3476_ _3526_ VGND VGND VPWR 
+ VPWR
+ _4320_ sky130_fd_sc_hd__a21oi_1
X_8701_ _3636_ _4320_ _3644_ _4150_ _4235_ VGND 
+ VGND
+ VPWR VPWR _4321_ sky130_fd_sc_hd__a2111o_2
X_8702_ _4319_ _4321_ VGND VGND VPWR VPWR 
+ _4322_
+ sky130_fd_sc_hd__nor2_1
X_8703_ _3453_ _4141_ _3694_ _4066_ VGND VGND 
+ VPWR
+ VPWR _4323_ sky130_fd_sc_hd__or4_1
X_8704_ _3703_ _4065_ VGND VGND VPWR VPWR 
+ _4324_
+ sky130_fd_sc_hd__or2_1
X_8705_ _3967_ _4230_ _4324_ _4165_ VGND VGND 
+ VPWR
+ VPWR _4325_ sky130_fd_sc_hd__or4_1
X_8706_ _4108_ _4242_ _4323_ _4325_ VGND VGND 
+ VPWR
+ VPWR _4326_ sky130_fd_sc_hd__or4_1
X_8707_ _4241_ _4229_ _4326_ VGND VGND VPWR 
+ VPWR
+ _4327_ sky130_fd_sc_hd__or3_2
X_8708_ _4020_ _3740_ _3684_ _3794_ VGND VGND 
+ VPWR
+ VPWR _4328_ sky130_fd_sc_hd__or4_1
X_8709_ _4180_ _4328_ _4254_ _4308_ VGND VGND 
+ VPWR
+ VPWR _4329_ sky130_fd_sc_hd__or4_1
X_8710_ _4247_ VGND VGND VPWR VPWR _4330_ sky130_fd_sc_hd__inv_2
X_8711_ _3630_ _4248_ _3746_ _4249_ _4330_ VGND 
+ VGND
+ VPWR VPWR _4331_ sky130_fd_sc_hd__o221ai_4
X_8712_ _4329_ _4331_ VGND VGND VPWR VPWR 
+ _4332_
+ sky130_fd_sc_hd__nor2_1
X_8713_ _3701_ _4187_ _4309_ _4186_ VGND VGND 
+ VPWR
+ VPWR _4333_ sky130_fd_sc_hd__or4_1
X_8714_ _4258_ _4333_ _4260_ _4310_ VGND VGND 
+ VPWR
+ VPWR _4334_ sky130_fd_sc_hd__or4_1
X_8715_ _3796_ _3902_ _3999_ VGND VGND VPWR 
+ VPWR
+ _4335_ sky130_fd_sc_hd__or3_1
X_8716_ _4205_ _4335_ _4269_ _4297_ VGND VGND 
+ VPWR
+ VPWR _4336_ sky130_fd_sc_hd__or4_1
X_8717_ _3738_ _3584_ _3738_ _3710_ VGND VGND 
+ VPWR
+ VPWR _4337_ sky130_fd_sc_hd__o22a_1
X_8718_ _3975_ _4337_ _3852_ _3841_ VGND VGND 
+ VPWR
+ VPWR _4338_ sky130_fd_sc_hd__o211ai_1
X_8719_ _4195_ _4338_ _4265_ VGND VGND VPWR 
+ VPWR
+ _4339_ sky130_fd_sc_hd__or3_2
X_8720_ _3724_ _4191_ _4006_ VGND VGND VPWR 
+ VPWR
+ _4340_ sky130_fd_sc_hd__or3_1
X_8721_ _3832_ _4211_ _4104_ _4340_ VGND VGND 
+ VPWR
+ VPWR _4341_ sky130_fd_sc_hd__or4_1
X_8722_ _3968_ _4274_ _4341_ VGND VGND VPWR 
+ VPWR
+ _4342_ sky130_fd_sc_hd__or3_1
X_8723_ _4303_ _4342_ _4300_ VGND VGND VPWR 
+ VPWR
+ _4343_ sky130_fd_sc_hd__nor3_4
X_8724_ _4336_ _4339_ _4343_ VGND VGND VPWR 
+ VPWR
+ _4344_ sky130_fd_sc_hd__o21ai_1
X_8725_ _4322_ _4327_ _4332_ _4334_ _4344_ VGND 
+ VGND
+ VPWR VPWR _0189_ sky130_fd_sc_hd__o221ai_1
X_8726_ _3478_ _3501_ _3872_ _3943_ _4130_ VGND 
+ VGND
+ VPWR VPWR _4345_ sky130_fd_sc_hd__o2111ai_4
X_8727_ _4221_ _4345_ _4282_ _4316_ VGND VGND 
+ VPWR
+ VPWR _4346_ sky130_fd_sc_hd__or4_1
X_8728_ _4346_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
X_8729_ _4336_ VGND VGND VPWR VPWR _4347_ sky130_fd_sc_hd__inv_2
X_8730_ _3769_ _3870_ _3989_ _4200_ VGND VGND 
+ VPWR
+ VPWR _4348_ sky130_fd_sc_hd__or4_2
X_8731_ _4266_ _4348_ _4339_ _4299_ VGND VGND 
+ VPWR
+ VPWR _4349_ sky130_fd_sc_hd__or4_1
X_8732_ _4319_ VGND VGND VPWR VPWR _4350_ sky130_fd_sc_hd__inv_2
X_8733_ _4327_ VGND VGND VPWR VPWR _4351_ sky130_fd_sc_hd__inv_2
X_8734_ _3502_ _4038_ _4084_ _4155_ VGND VGND 
+ VPWR
+ VPWR _4352_ sky130_fd_sc_hd__or4_1
X_8735_ _4231_ _4352_ _4321_ _4288_ VGND VGND 
+ VPWR
+ VPWR _4353_ sky130_fd_sc_hd__or4_1
X_8736_ _3584_ _3621_ _3659_ _4039_ VGND VGND 
+ VPWR
+ VPWR _4354_ sky130_fd_sc_hd__o211a_1
X_8737_ _3623_ _4171_ _4354_ _4252_ VGND VGND 
+ VPWR
+ VPWR _4355_ sky130_fd_sc_hd__o211ai_4
X_8738_ _4329_ VGND VGND VPWR VPWR _4356_ sky130_fd_sc_hd__inv_2
X_8739_ _4334_ VGND VGND VPWR VPWR _4357_ sky130_fd_sc_hd__inv_2
X_8740_ _4331_ _4355_ _4306_ _4356_ _4357_ VGND 
+ VGND
+ VPWR VPWR _4358_ sky130_fd_sc_hd__o311a_1
X_8741_ _4350_ _4351_ _4353_ _4358_ VGND VGND 
+ VPWR
+ VPWR _4359_ sky130_fd_sc_hd__a31o_1
X_8742_ _4347_ _4343_ _4349_ _4359_ VGND VGND 
+ VPWR
+ VPWR _0191_ sky130_fd_sc_hd__a31o_1
X_8743_ _4408_ VGND VGND VPWR VPWR _4360_ sky130_fd_sc_hd__clkbuf_1
X_8744_ _4360_ VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__clkbuf_1
X_8745_ _4411_ VGND VGND VPWR VPWR _4361_ sky130_fd_sc_hd__clkbuf_1
X_8746_ _4361_ VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__clkbuf_1
X_8747_ _4414_ VGND VGND VPWR VPWR _4362_ sky130_fd_sc_hd__clkbuf_1
X_8748_ _4362_ VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__clkbuf_1
X_8749_ _4415_ VGND VGND VPWR VPWR _4363_ sky130_fd_sc_hd__clkbuf_1
X_8750_ _4363_ VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__clkbuf_1
X_8751_ _4416_ VGND VGND VPWR VPWR _4364_ sky130_fd_sc_hd__clkbuf_1
X_8752_ _4364_ VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__clkbuf_1
X_8753_ _4417_ VGND VGND VPWR VPWR _4365_ sky130_fd_sc_hd__clkbuf_1
X_8754_ _4365_ VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__clkbuf_1
X_8755_ _4418_ VGND VGND VPWR VPWR _4366_ sky130_fd_sc_hd__clkbuf_1
X_8756_ _4366_ VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__clkbuf_1
X_8757_ _4419_ VGND VGND VPWR VPWR _4367_ sky130_fd_sc_hd__clkbuf_1
X_8758_ _4367_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__clkbuf_1
X_8759_ _4420_ VGND VGND VPWR VPWR _4368_ sky130_fd_sc_hd__clkbuf_1
X_8760_ _4368_ VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__clkbuf_1
X_8761_ _4421_ VGND VGND VPWR VPWR _4369_ sky130_fd_sc_hd__clkbuf_1
X_8762_ _4369_ VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__clkbuf_1
X_8763_ _4422_ VGND VGND VPWR VPWR _4370_ sky130_fd_sc_hd__clkbuf_1
X_8764_ _4370_ VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__clkbuf_1
X_8765_ _4423_ VGND VGND VPWR VPWR _4371_ sky130_fd_sc_hd__clkbuf_1
X_8766_ _4371_ VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__clkbuf_1
X_8767_ _4424_ VGND VGND VPWR VPWR _4372_ sky130_fd_sc_hd__clkbuf_1
X_8768_ _4372_ VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__clkbuf_1
X_8769_ _4425_ VGND VGND VPWR VPWR _4373_ sky130_fd_sc_hd__clkbuf_1
X_8770_ _4373_ VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__clkbuf_1
X_8771_ _4426_ VGND VGND VPWR VPWR _4374_ sky130_fd_sc_hd__clkbuf_1
X_8772_ _4374_ VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__clkbuf_1
X_8773_ _4427_ VGND VGND VPWR VPWR _4375_ sky130_fd_sc_hd__clkbuf_1
X_8774_ _4375_ VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__clkbuf_1
X_8775_ _4428_ VGND VGND VPWR VPWR _4376_ sky130_fd_sc_hd__clkbuf_1
X_8776_ _4376_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__clkbuf_1
X_8777_ _4429_ VGND VGND VPWR VPWR _4377_ sky130_fd_sc_hd__clkbuf_1
X_8778_ _4377_ VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__clkbuf_1
X_8779_ _4430_ VGND VGND VPWR VPWR _4378_ sky130_fd_sc_hd__clkbuf_1
X_8780_ _4378_ VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__clkbuf_1
X_8781_ _4431_ VGND VGND VPWR VPWR _4379_ sky130_fd_sc_hd__clkbuf_1
X_8782_ _4379_ VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__clkbuf_1
X_8783_ _4432_ VGND VGND VPWR VPWR _4380_ sky130_fd_sc_hd__clkbuf_1
X_8784_ _4380_ VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__clkbuf_1
X_8785_ _4433_ VGND VGND VPWR VPWR _4381_ sky130_fd_sc_hd__clkbuf_1
X_8786_ _4381_ VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__clkbuf_1
X_8787_ _4434_ VGND VGND VPWR VPWR _4382_ sky130_fd_sc_hd__clkbuf_1
X_8788_ _4382_ VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__clkbuf_1
X_8789_ _4435_ VGND VGND VPWR VPWR _4383_ sky130_fd_sc_hd__clkbuf_1
X_8790_ _4383_ VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__clkbuf_1
X_8791_ _4436_ VGND VGND VPWR VPWR _4384_ sky130_fd_sc_hd__clkbuf_1
X_8792_ _4384_ VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__clkbuf_1
X_8793_ _4437_ VGND VGND VPWR VPWR _4385_ sky130_fd_sc_hd__clkbuf_1
X_8794_ _4385_ VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__clkbuf_1
X_8795_ _4438_ VGND VGND VPWR VPWR _4386_ sky130_fd_sc_hd__clkbuf_1
X_8796_ _4386_ VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__clkbuf_1
X_8797_ _4439_ VGND VGND VPWR VPWR _4387_ sky130_fd_sc_hd__clkbuf_1
X_8798_ _4387_ VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__clkbuf_1
X_8799_ _4440_ VGND VGND VPWR VPWR _4388_ sky130_fd_sc_hd__clkbuf_1
X_8800_ _4388_ VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__clkbuf_1
X_8801_ net68 net126 VGND VGND VPWR VPWR 
+ _4389_
+ sky130_fd_sc_hd__and2_1
X_8802_ _4389_ VGND VGND VPWR VPWR net305 sky130_fd_sc_hd__clkbuf_1
X_8803_ net63 net79 VGND VGND VPWR VPWR 
+ _4390_
+ sky130_fd_sc_hd__and2_1
X_8804_ _4390_ VGND VGND VPWR VPWR net311 sky130_fd_sc_hd__clkbuf_1
X_8805_ net36 net1 VGND VGND VPWR VPWR 
+ _4391_
+ sky130_fd_sc_hd__and2_1
X_8806_ _4391_ VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__clkbuf_1
X_8807_ _1303_ _1848_ VGND VGND VPWR VPWR 
+ net205
+ sky130_fd_sc_hd__nor2_2
X_8808_ _2597_ _2233_ VGND VGND VPWR VPWR 
+ net206
+ sky130_fd_sc_hd__nor2_2
X_8809_ _2693_ VGND VGND VPWR VPWR _4392_ sky130_fd_sc_hd__inv_2
X_8810_ _1082_ _4392_ VGND VGND VPWR VPWR 
+ _0027_
+ sky130_fd_sc_hd__nor2_1
X_8811_ _1081_ _4392_ VGND VGND VPWR VPWR 
+ _0026_
+ sky130_fd_sc_hd__nor2_1
X_8812_ _1083_ _4392_ VGND VGND VPWR VPWR 
+ _0025_
+ sky130_fd_sc_hd__nor2_1
X_8813_ _1084_ _4392_ VGND VGND VPWR VPWR 
+ _0024_
+ sky130_fd_sc_hd__nor2_1
X_8814_ serial_xfer _2032_ net368 _1032_ _0063_ VGND 
+ VGND
+ VPWR VPWR _1020_ sky130_fd_sc_hd__o221a_1
X_8815__378 VGND VGND VPWR VPWR net378 NC sky130_fd_sc_hd__conb_1
X_8816_ net87 VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__clkbuf_1
X_8817_ net65 VGND VGND VPWR VPWR net314 sky130_fd_sc_hd__clkbuf_1
X_8818_ net66 VGND VGND VPWR VPWR net315 sky130_fd_sc_hd__clkbuf_1
X_8819_ serial_clock_pre serial_bb_clock serial_bb_enable VGND VGND VPWR 
+ VPWR
+ net306 sky130_fd_sc_hd__mux2_1
X_8820_ serial_load_pre serial_bb_load serial_bb_enable VGND VGND VPWR 
+ VPWR
+ net309 sky130_fd_sc_hd__mux2_1
X_8821_ serial_resetn_pre serial_bb_resetn serial_bb_enable VGND VGND VPWR 
+ VPWR
+ net310 sky130_fd_sc_hd__mux2_1
X_8822_ \serial_data_staging_1[12]\ serial_bb_data_1 serial_bb_enable VGND VGND VPWR 
+ VPWR
+ net307 sky130_fd_sc_hd__mux2_4
X_8823_ \serial_data_staging_2[12]\ serial_bb_data_2 serial_bb_enable VGND VGND VPWR 
+ VPWR
+ net308 sky130_fd_sc_hd__mux2_1
X_8824_ \mgmt_gpio_data[0]\ net3 net1 VGND VGND VPWR 
+ VPWR
+ net245 sky130_fd_sc_hd__mux2_2
X_8825_ \mgmt_gpio_data[1]\ \hkspi.SDO\ _0079_ VGND VGND VPWR 
+ VPWR
+ _0095_ sky130_fd_sc_hd__mux2_1
X_8826_ _0095_ net38 \hkspi.pass_thru_user\ VGND VGND VPWR 
+ VPWR
+ _0096_ sky130_fd_sc_hd__mux2_1
X_8827_ _0096_ net74 \hkspi.pass_thru_mgmt\ VGND VGND VPWR 
+ VPWR
+ net246 sky130_fd_sc_hd__mux2_4
X_8828_ \mgmt_gpio_data[35]\ net81 net79 VGND VGND VPWR 
+ VPWR
+ net247 sky130_fd_sc_hd__mux2_1
X_8829_ \mgmt_gpio_data[36]\ net89 net76 VGND VGND VPWR 
+ VPWR
+ net248 sky130_fd_sc_hd__mux2_1
X_8830_ \mgmt_gpio_data[37]\ net91 net76 VGND VGND VPWR 
+ VPWR
+ net249 sky130_fd_sc_hd__mux2_1
X_8831_ _0097_ net2 net1 VGND VGND VPWR 
+ VPWR
+ net207 sky130_fd_sc_hd__mux2_2
X_8832_ _0097_ \hkspi.sdoenb\ _0079_ VGND VGND VPWR 
+ VPWR
+ net218 sky130_fd_sc_hd__mux2_1
X_8833_ _0094_ net82 net79 VGND VGND VPWR 
+ VPWR
+ net235 sky130_fd_sc_hd__mux2_4
X_8834_ _0093_ net90 net76 VGND VGND VPWR 
+ VPWR
+ net236 sky130_fd_sc_hd__mux2_2
X_8835_ _0092_ net92 net76 VGND VGND VPWR 
+ VPWR
+ net237 sky130_fd_sc_hd__mux2_1
X_8836_ net84 net67 \hkspi.pass_thru_mgmt_delay\ VGND VGND VPWR 
+ VPWR
+ net252 sky130_fd_sc_hd__mux2_2
X_8837_ net83 clknet_2_0_0_mgmt_gpio_in[4] \hkspi.pass_thru_mgmt\ VGND VGND VPWR 
+ VPWR
+ net250 sky130_fd_sc_hd__mux2_1
X_8838_ net85 net58 \hkspi.pass_thru_mgmt_delay\ VGND VGND VPWR 
+ VPWR
+ net254 sky130_fd_sc_hd__mux2_2
X_8839_ net58 \wbbd_data[0]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[0]\ sky130_fd_sc_hd__mux2_8
X_8840_ \hkspi.odata[1]\ \wbbd_data[1]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[1]\ sky130_fd_sc_hd__mux2_8
X_8841_ \hkspi.odata[2]\ \wbbd_data[2]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[2]\ sky130_fd_sc_hd__mux2_8
X_8842_ \hkspi.odata[3]\ \wbbd_data[3]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[3]\ sky130_fd_sc_hd__mux2_8
X_8843_ \hkspi.odata[4]\ \wbbd_data[4]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[4]\ sky130_fd_sc_hd__mux2_8
X_8844_ \hkspi.odata[5]\ \wbbd_data[5]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[5]\ sky130_fd_sc_hd__mux2_8
X_8845_ \hkspi.odata[6]\ \wbbd_data[6]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[6]\ sky130_fd_sc_hd__mux2_8
X_8846_ \hkspi.odata[7]\ \wbbd_data[7]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ \cdata[7]\ sky130_fd_sc_hd__mux2_8
X_8847_ _0098_ wbbd_sck wbbd_busy VGND VGND VPWR 
+ VPWR
+ csclk sky130_fd_sc_hd__mux2_1
X_8848_ \mgmt_gpio_data_buf[16]\ net368 _0080_ VGND VGND VPWR 
+ VPWR
+ _0208_ sky130_fd_sc_hd__mux2_1
X_8849_ \mgmt_gpio_data_buf[0]\ net368 _0085_ VGND VGND VPWR 
+ VPWR
+ _0192_ sky130_fd_sc_hd__mux2_1
X_8850_ _0130_ \gpio_configure[0][1]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0131_ sky130_fd_sc_hd__mux2_1
X_8851_ _0131_ \serial_data_staging_1[0]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0003_ sky130_fd_sc_hd__mux2_1
X_8852_ _0132_ \gpio_configure[0][2]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0133_ sky130_fd_sc_hd__mux2_1
X_8853_ _0133_ \serial_data_staging_1[1]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0004_ sky130_fd_sc_hd__mux2_1
X_8854_ _0134_ \gpio_configure[0][3]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0135_ sky130_fd_sc_hd__mux2_1
X_8855_ _0135_ \serial_data_staging_1[2]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0005_ sky130_fd_sc_hd__mux2_1
X_8856_ _0136_ \gpio_configure[0][4]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0137_ sky130_fd_sc_hd__mux2_1
X_8857_ _0137_ \serial_data_staging_1[3]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0006_ sky130_fd_sc_hd__mux2_1
X_8858_ _0138_ \gpio_configure[0][5]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0139_ sky130_fd_sc_hd__mux2_1
X_8859_ _0139_ \serial_data_staging_1[4]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0007_ sky130_fd_sc_hd__mux2_1
X_8860_ _0140_ \gpio_configure[0][6]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0141_ sky130_fd_sc_hd__mux2_1
X_8861_ _0141_ \serial_data_staging_1[5]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0008_ sky130_fd_sc_hd__mux2_1
X_8862_ _0142_ \gpio_configure[0][7]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0143_ sky130_fd_sc_hd__mux2_1
X_8863_ _0143_ \serial_data_staging_1[6]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0009_ sky130_fd_sc_hd__mux2_1
X_8864_ _0144_ \gpio_configure[0][8]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0145_ sky130_fd_sc_hd__mux2_1
X_8865_ _0145_ \serial_data_staging_1[7]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0010_ sky130_fd_sc_hd__mux2_1
X_8866_ _0146_ \gpio_configure[0][9]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0147_ sky130_fd_sc_hd__mux2_1
X_8867_ _0147_ \serial_data_staging_1[8]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0011_ sky130_fd_sc_hd__mux2_1
X_8868_ _0148_ \gpio_configure[0][10]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0149_ sky130_fd_sc_hd__mux2_1
X_8869_ _0149_ \serial_data_staging_1[9]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0000_ sky130_fd_sc_hd__mux2_1
X_8870_ _0150_ \gpio_configure[0][11]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0151_ sky130_fd_sc_hd__mux2_1
X_8871_ _0151_ \serial_data_staging_1[10]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0001_ sky130_fd_sc_hd__mux2_1
X_8872_ _0152_ \gpio_configure[0][12]\ _0127_ VGND VGND VPWR 
+ VPWR
+ _0153_ sky130_fd_sc_hd__mux2_1
X_8873_ _0153_ \serial_data_staging_1[11]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0002_ sky130_fd_sc_hd__mux2_1
X_8874_ _0103_ \gpio_configure[0][1]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0104_ sky130_fd_sc_hd__mux2_1
X_8875_ _0104_ \serial_data_staging_2[0]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0015_ sky130_fd_sc_hd__mux2_1
X_8876_ _0105_ \gpio_configure[0][2]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0106_ sky130_fd_sc_hd__mux2_1
X_8877_ _0106_ \serial_data_staging_2[1]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0016_ sky130_fd_sc_hd__mux2_1
X_8878_ _0107_ \gpio_configure[0][3]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0108_ sky130_fd_sc_hd__mux2_1
X_8879_ _0108_ \serial_data_staging_2[2]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0017_ sky130_fd_sc_hd__mux2_1
X_8880_ _0109_ \gpio_configure[0][4]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0110_ sky130_fd_sc_hd__mux2_1
X_8881_ _0110_ \serial_data_staging_2[3]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0018_ sky130_fd_sc_hd__mux2_1
X_8882_ _0111_ \gpio_configure[0][5]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0112_ sky130_fd_sc_hd__mux2_1
X_8883_ _0112_ \serial_data_staging_2[4]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0019_ sky130_fd_sc_hd__mux2_1
X_8884_ _0113_ \gpio_configure[0][6]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0114_ sky130_fd_sc_hd__mux2_1
X_8885_ _0114_ \serial_data_staging_2[5]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0020_ sky130_fd_sc_hd__mux2_1
X_8886_ _0115_ \gpio_configure[0][7]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0116_ sky130_fd_sc_hd__mux2_1
X_8887_ _0116_ \serial_data_staging_2[6]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0021_ sky130_fd_sc_hd__mux2_1
X_8888_ _0117_ \gpio_configure[0][8]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0118_ sky130_fd_sc_hd__mux2_1
X_8889_ _0118_ \serial_data_staging_2[7]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0022_ sky130_fd_sc_hd__mux2_1
X_8890_ _0119_ \gpio_configure[0][9]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0120_ sky130_fd_sc_hd__mux2_1
X_8891_ _0120_ \serial_data_staging_2[8]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0023_ sky130_fd_sc_hd__mux2_1
X_8892_ _0121_ \gpio_configure[0][10]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0122_ sky130_fd_sc_hd__mux2_1
X_8893_ _0122_ \serial_data_staging_2[9]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0012_ sky130_fd_sc_hd__mux2_1
X_8894_ _0123_ \gpio_configure[0][11]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0124_ sky130_fd_sc_hd__mux2_1
X_8895_ _0124_ \serial_data_staging_2[10]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0013_ sky130_fd_sc_hd__mux2_1
X_8896_ _0125_ \gpio_configure[0][12]\ _0100_ VGND VGND VPWR 
+ VPWR
+ _0126_ sky130_fd_sc_hd__mux2_1
X_8897_ _0126_ \serial_data_staging_2[11]\ \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0014_ sky130_fd_sc_hd__mux2_1
X_8898_ \mgmt_gpio_data_buf[15]\ \cdata[7]\ _0083_ VGND VGND VPWR 
+ VPWR
+ _0207_ sky130_fd_sc_hd__mux2_1
X_8899_ _0158_ \hkspi.addr[1]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0049_ sky130_fd_sc_hd__mux2_1
X_8900_ _0157_ \hkspi.addr[0]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0048_ sky130_fd_sc_hd__mux2_1
X_8901_ _0165_ \hkspi.fixed[0]\ \hkspi.state[0]\ VGND VGND VPWR 
+ VPWR
+ _0044_ sky130_fd_sc_hd__mux2_1
X_8902_ _0156_ net58 \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0047_ sky130_fd_sc_hd__mux2_1
X_8903_ \mgmt_gpio_data_buf[1]\ net366 _0085_ VGND VGND VPWR 
+ VPWR
+ _0193_ sky130_fd_sc_hd__mux2_1
X_8904_ \mgmt_gpio_data_buf[6]\ \cdata[6]\ _0085_ VGND VGND VPWR 
+ VPWR
+ _0198_ sky130_fd_sc_hd__mux2_1
X_8905_ \mgmt_gpio_data_buf[10]\ net364 _0083_ VGND VGND VPWR 
+ VPWR
+ _0202_ sky130_fd_sc_hd__mux2_1
X_8906_ \mgmt_gpio_data_buf[12]\ net360 _0083_ VGND VGND VPWR 
+ VPWR
+ _0204_ sky130_fd_sc_hd__mux2_1
X_8907_ _0163_ \hkspi.addr[6]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0054_ sky130_fd_sc_hd__mux2_1
X_8908_ _0164_ net58 \hkspi.state[0]\ VGND VGND VPWR 
+ VPWR
+ _0043_ sky130_fd_sc_hd__mux2_1
X_8909_ _0166_ \hkspi.fixed[1]\ \hkspi.state[0]\ VGND VGND VPWR 
+ VPWR
+ _0045_ sky130_fd_sc_hd__mux2_1
X_8910_ _0159_ \hkspi.addr[2]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0050_ sky130_fd_sc_hd__mux2_1
X_8911_ _0160_ \hkspi.addr[3]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0051_ sky130_fd_sc_hd__mux2_1
X_8912_ _0161_ \hkspi.addr[4]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0052_ sky130_fd_sc_hd__mux2_1
X_8913_ _0162_ \hkspi.addr[5]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0053_ sky130_fd_sc_hd__mux2_1
X_8914_ \mgmt_gpio_data_buf[7]\ \cdata[7]\ _0085_ VGND VGND VPWR 
+ VPWR
+ _0199_ sky130_fd_sc_hd__mux2_1
X_8915_ \mgmt_gpio_data_buf[5]\ \cdata[5]\ _0085_ VGND VGND VPWR 
+ VPWR
+ _0197_ sky130_fd_sc_hd__mux2_1
X_8916_ \mgmt_gpio_data_buf[8]\ net368 _0083_ VGND VGND VPWR 
+ VPWR
+ _0200_ sky130_fd_sc_hd__mux2_1
X_8917_ \mgmt_gpio_data_buf[23]\ \cdata[7]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0215_ sky130_fd_sc_hd__mux2_1
X_8918_ \mgmt_gpio_data_buf[22]\ \cdata[6]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0214_ sky130_fd_sc_hd__mux2_1
X_8919_ \mgmt_gpio_data_buf[17]\ \cdata[1]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0209_ sky130_fd_sc_hd__mux2_1
X_8920_ \mgmt_gpio_data_buf[4]\ net360 _0085_ VGND VGND VPWR 
+ VPWR
+ _0196_ sky130_fd_sc_hd__mux2_1
X_8921_ \mgmt_gpio_data_buf[21]\ \cdata[5]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0213_ sky130_fd_sc_hd__mux2_1
X_8922_ \mgmt_gpio_data_buf[18]\ \cdata[2]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0210_ sky130_fd_sc_hd__mux2_1
X_8923_ \mgmt_gpio_data_buf[3]\ net362 _0085_ VGND VGND VPWR 
+ VPWR
+ _0195_ sky130_fd_sc_hd__mux2_1
X_8924_ \xfer_state[2]\ net306 \xfer_state[1]\ VGND VGND VPWR 
+ VPWR
+ _0042_ sky130_fd_sc_hd__mux2_1
X_8925_ \mgmt_gpio_data_buf[20]\ net360 _0080_ VGND VGND VPWR 
+ VPWR
+ _0212_ sky130_fd_sc_hd__mux2_1
X_8926_ \mgmt_gpio_data_buf[19]\ \cdata[3]\ _0080_ VGND VGND VPWR 
+ VPWR
+ _0211_ sky130_fd_sc_hd__mux2_1
X_8927_ \mgmt_gpio_data_buf[14]\ \cdata[6]\ _0083_ VGND VGND VPWR 
+ VPWR
+ _0206_ sky130_fd_sc_hd__mux2_1
X_8928_ \mgmt_gpio_data_buf[13]\ \cdata[5]\ _0083_ VGND VGND VPWR 
+ VPWR
+ _0205_ sky130_fd_sc_hd__mux2_1
X_8929_ \mgmt_gpio_data_buf[11]\ net362 _0083_ VGND VGND VPWR 
+ VPWR
+ _0203_ sky130_fd_sc_hd__mux2_1
X_8930_ \mgmt_gpio_data_buf[9]\ net366 _0083_ VGND VGND VPWR 
+ VPWR
+ _0201_ sky130_fd_sc_hd__mux2_1
X_8931_ \hkspi.addr[2]\ \hkspi.addr[1]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0068_ sky130_fd_sc_hd__mux2_1
X_8932_ _0068_ \wbbd_addr[2]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0069_ sky130_fd_sc_hd__mux2_4
X_8933_ \hkspi.addr[3]\ \hkspi.addr[2]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0070_ sky130_fd_sc_hd__mux2_1
X_8934_ _0070_ \wbbd_addr[3]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0071_ sky130_fd_sc_hd__mux2_4
X_8935_ \hkspi.addr[4]\ \hkspi.addr[3]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0072_ sky130_fd_sc_hd__mux2_1
X_8936_ _0072_ \wbbd_addr[4]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0073_ sky130_fd_sc_hd__mux2_2
X_8937_ \hkspi.addr[5]\ \hkspi.addr[4]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0074_ sky130_fd_sc_hd__mux2_1
X_8938_ _0074_ \wbbd_addr[5]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0075_ sky130_fd_sc_hd__mux2_2
X_8939_ \hkspi.wrstb\ wbbd_write wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0063_ sky130_fd_sc_hd__mux2_8
X_8940_ \hkspi.addr[6]\ \hkspi.addr[5]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0076_ sky130_fd_sc_hd__mux2_1
X_8941_ _0076_ \wbbd_addr[6]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0077_ sky130_fd_sc_hd__mux2_1
X_8942_ \hkspi.addr[7]\ \hkspi.addr[6]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0078_ sky130_fd_sc_hd__mux2_1
X_8943_ \hkspi.addr[0]\ net58 \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0064_ sky130_fd_sc_hd__mux2_1
X_8944_ _0064_ \wbbd_addr[0]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0065_ sky130_fd_sc_hd__mux2_4
X_8945_ \hkspi.addr[1]\ \hkspi.addr[0]\ \hkspi.state[3]\ VGND VGND VPWR 
+ VPWR
+ _0066_ sky130_fd_sc_hd__mux2_1
X_8946_ _0066_ \wbbd_addr[1]\ wbbd_busy VGND VGND VPWR 
+ VPWR
+ _0067_ sky130_fd_sc_hd__mux2_4
X_8947_ \hkspi.ldata[4]\ \hkspi.idata[5]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0059_ sky130_fd_sc_hd__mux2_1
X_8948_ net393 \hkspi.idata[6]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0060_ sky130_fd_sc_hd__mux2_1
X_8949_ \hkspi.ldata[2]\ \hkspi.idata[3]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0057_ sky130_fd_sc_hd__mux2_1
X_8950_ \hkspi.ldata[3]\ \hkspi.idata[4]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0058_ sky130_fd_sc_hd__mux2_1
X_8951_ \hkspi.ldata[1]\ \hkspi.idata[2]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0056_ sky130_fd_sc_hd__mux2_1
X_8952_ \hkspi.ldata[0]\ \hkspi.idata[1]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0055_ sky130_fd_sc_hd__mux2_1
X_8953_ \hkspi.ldata[6]\ \hkspi.idata[7]\ _0062_ VGND VGND VPWR 
+ VPWR
+ _0061_ sky130_fd_sc_hd__mux2_1
X_8954_ _0155_ _0154_ \hkspi.state[2]\ VGND VGND VPWR 
+ VPWR
+ _0046_ sky130_fd_sc_hd__mux2_1
X_8955_ \mgmt_gpio_data_buf[2]\ net364 _0085_ VGND VGND VPWR 
+ VPWR
+ _0194_ sky130_fd_sc_hd__mux2_1
X_8956_ _0085_ _0081_ _0079_ VGND VGND VPWR 
+ VPWR
+ _0086_ sky130_fd_sc_hd__mux2_1
X_8957_ _0089_ _0087_ _0062_ VGND VGND VPWR 
+ VPWR
+ _0090_ sky130_fd_sc_hd__mux2_1
X_8958_ \hkspi.count[0]\ \hkspi.count[2]\ \hkspi.count[1]\ VGND VGND VPWR 
+ VPWR
+ _0091_ sky130_fd_sc_hd__mux2_1
X_8959_ _0101_ _0099_ _0100_ VGND VGND VPWR 
+ VPWR
+ _0102_ sky130_fd_sc_hd__mux2_1
X_8960_ _0168_ _0088_ _0167_ VGND VGND VPWR 
+ VPWR
+ _4442_ sky130_fd_sc_hd__mux2_1
X_8961_ _0170_ net164 _0169_ VGND VGND VPWR 
+ VPWR
+ _4393_ sky130_fd_sc_hd__mux2_1
X_8962_ _0171_ net175 _0169_ VGND VGND VPWR 
+ VPWR
+ _4394_ sky130_fd_sc_hd__mux2_1
X_8963_ _0172_ net186 _0169_ VGND VGND VPWR 
+ VPWR
+ _4395_ sky130_fd_sc_hd__mux2_1
X_8964_ _0173_ net189 _0169_ VGND VGND VPWR 
+ VPWR
+ _4396_ sky130_fd_sc_hd__mux2_1
X_8965_ _0174_ net190 _0169_ VGND VGND VPWR 
+ VPWR
+ _4397_ sky130_fd_sc_hd__mux2_1
X_8966_ _0175_ net191 _0169_ VGND VGND VPWR 
+ VPWR
+ _4398_ sky130_fd_sc_hd__mux2_1
X_8967_ _0176_ net192 _0169_ VGND VGND VPWR 
+ VPWR
+ _4399_ sky130_fd_sc_hd__mux2_1
X_8968_ _0177_ net193 _0169_ VGND VGND VPWR 
+ VPWR
+ _4400_ sky130_fd_sc_hd__mux2_1
X_8969_ _0179_ _0178_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4401_ sky130_fd_sc_hd__mux2_4
X_8970_ _0181_ _0180_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4402_ sky130_fd_sc_hd__mux2_4
X_8971_ _0183_ _0182_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4403_ sky130_fd_sc_hd__mux2_4
X_8972_ _0185_ _0184_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4404_ sky130_fd_sc_hd__mux2_2
X_8973_ _0187_ _0186_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4405_ sky130_fd_sc_hd__mux2_2
X_8974_ _0189_ _0188_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4406_ sky130_fd_sc_hd__mux2_2
X_8975_ _0191_ _0190_ _0169_ VGND VGND VPWR 
+ VPWR
+ _4407_ sky130_fd_sc_hd__mux2_2
X_8976_ _0080_ _0081_ _0079_ VGND VGND VPWR 
+ VPWR
+ _0082_ sky130_fd_sc_hd__mux2_1
X_8977_ _0083_ _0081_ _0079_ VGND VGND VPWR 
+ VPWR
+ _0084_ sky130_fd_sc_hd__mux2_1
X_8978_ _0128_ _0099_ _0127_ VGND VGND VPWR 
+ VPWR
+ _0129_ sky130_fd_sc_hd__mux2_1
X_8979_ \mgmt_gpio_data[2]\ _4408_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[2]
+ sky130_fd_sc_hd__ebufn_8
X_8980_ \mgmt_gpio_data[3]\ _4409_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[3]
+ sky130_fd_sc_hd__ebufn_8
X_8981_ \mgmt_gpio_data[4]\ _4410_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[4]
+ sky130_fd_sc_hd__ebufn_8
X_8982_ \mgmt_gpio_data[5]\ _4411_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[5]
+ sky130_fd_sc_hd__ebufn_8
X_8983_ \mgmt_gpio_out_pre[6]\ _4412_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[6]
+ sky130_fd_sc_hd__ebufn_8
X_8984_ \mgmt_gpio_data[7]\ _4413_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[7]
+ sky130_fd_sc_hd__ebufn_8
X_8985_ \mgmt_gpio_out_pre[8]\ _4414_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[8]
+ sky130_fd_sc_hd__ebufn_8
X_8986_ \mgmt_gpio_out_pre[9]\ _4415_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[9]
+ sky130_fd_sc_hd__ebufn_2
X_8987_ \mgmt_gpio_out_pre[10]\ _4416_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[10]
+ sky130_fd_sc_hd__ebufn_8
X_8988_ \mgmt_gpio_data[11]\ _4417_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[11]
+ sky130_fd_sc_hd__ebufn_8
X_8989_ \mgmt_gpio_data[12]\ _4418_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[12]
+ sky130_fd_sc_hd__ebufn_8
X_8990_ \mgmt_gpio_out_pre[13]\ _4419_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[13]
+ sky130_fd_sc_hd__ebufn_8
X_8991_ \mgmt_gpio_out_pre[14]\ _4420_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[14]
+ sky130_fd_sc_hd__ebufn_2
X_8992_ \mgmt_gpio_out_pre[15]\ _4421_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[15]
+ sky130_fd_sc_hd__ebufn_2
X_8993_ \mgmt_gpio_data[16]\ _4422_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[16]
+ sky130_fd_sc_hd__ebufn_8
X_8994_ \mgmt_gpio_data[17]\ _4423_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[17]
+ sky130_fd_sc_hd__ebufn_8
X_8995_ \mgmt_gpio_data[18]\ _4424_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[18]
+ sky130_fd_sc_hd__ebufn_8
X_8996_ \mgmt_gpio_data[19]\ _4425_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[19]
+ sky130_fd_sc_hd__ebufn_8
X_8997_ \mgmt_gpio_data[20]\ _4426_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[20]
+ sky130_fd_sc_hd__ebufn_8
X_8998_ \mgmt_gpio_data[21]\ _4427_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[21]
+ sky130_fd_sc_hd__ebufn_8
X_8999_ \mgmt_gpio_data[22]\ _4428_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[22]
+ sky130_fd_sc_hd__ebufn_8
X_9000_ \mgmt_gpio_data[23]\ _4429_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[23]
+ sky130_fd_sc_hd__ebufn_8
X_9001_ \mgmt_gpio_data[24]\ _4430_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[24]
+ sky130_fd_sc_hd__ebufn_8
X_9002_ \mgmt_gpio_data[25]\ _4431_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[25]
+ sky130_fd_sc_hd__ebufn_8
X_9003_ \mgmt_gpio_data[26]\ _4432_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[26]
+ sky130_fd_sc_hd__ebufn_8
X_9004_ \mgmt_gpio_data[27]\ _4433_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[27]
+ sky130_fd_sc_hd__ebufn_8
X_9005_ \mgmt_gpio_data[28]\ _4434_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[28]
+ sky130_fd_sc_hd__ebufn_8
X_9006_ \mgmt_gpio_data[29]\ _4435_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[29]
+ sky130_fd_sc_hd__ebufn_8
X_9007_ \mgmt_gpio_data[30]\ _4436_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[30]
+ sky130_fd_sc_hd__ebufn_8
X_9008_ \mgmt_gpio_data[31]\ _4437_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[31]
+ sky130_fd_sc_hd__ebufn_8
X_9009_ \mgmt_gpio_out_pre[32]\ _4438_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[32]
+ sky130_fd_sc_hd__ebufn_8
X_9010_ \mgmt_gpio_out_pre[33]\ _4439_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[33]
+ sky130_fd_sc_hd__ebufn_8
X_9011_ \mgmt_gpio_data[34]\ _4440_ VGND VGND VPWR VPWR 
+ mgmt_gpio_out[34]
+ sky130_fd_sc_hd__ebufn_8
X_9012_ clknet_3_4_0_wb_clk_i _0262_ VGND VGND VPWR VPWR 
+ net357
+ sky130_fd_sc_hd__dfxtp_1
X_9013_ clknet_3_5_0_wb_clk_i _0263_ VGND VGND VPWR VPWR 
+ net358
+ sky130_fd_sc_hd__dfxtp_1
X_9014_ clknet_3_4_0_wb_clk_i _0264_ VGND VGND VPWR VPWR 
+ net328
+ sky130_fd_sc_hd__dfxtp_1
X_9015_ clknet_3_5_0_wb_clk_i _0265_ VGND VGND VPWR VPWR 
+ net329
+ sky130_fd_sc_hd__dfxtp_1
X_9016_ clknet_3_5_0_wb_clk_i _0266_ VGND VGND VPWR VPWR 
+ net330
+ sky130_fd_sc_hd__dfxtp_1
X_9017_ clknet_3_7_0_wb_clk_i _0267_ VGND VGND VPWR VPWR 
+ net331
+ sky130_fd_sc_hd__dfxtp_1
X_9018_ clknet_3_5_0_wb_clk_i _0268_ VGND VGND VPWR VPWR 
+ net332
+ sky130_fd_sc_hd__dfxtp_1
X_9019_ clknet_3_5_0_wb_clk_i _0269_ VGND VGND VPWR VPWR 
+ net333
+ sky130_fd_sc_hd__dfxtp_1
X_9020_ clknet_3_4_0_wb_clk_i _0270_ VGND VGND VPWR VPWR 
+ net327
+ sky130_fd_sc_hd__dfxtp_1
X_9021_ clknet_3_4_0_wb_clk_i _0271_ VGND VGND VPWR VPWR 
+ net338
+ sky130_fd_sc_hd__dfxtp_1
X_9022_ clknet_3_4_0_wb_clk_i _0272_ VGND VGND VPWR VPWR 
+ net349
+ sky130_fd_sc_hd__dfxtp_1
X_9023_ clknet_3_4_0_wb_clk_i _0273_ VGND VGND VPWR VPWR 
+ net352
+ sky130_fd_sc_hd__dfxtp_1
X_9024_ clknet_3_4_0_wb_clk_i _0274_ VGND VGND VPWR VPWR 
+ net353
+ sky130_fd_sc_hd__dfxtp_1
X_9025_ clknet_3_4_0_wb_clk_i _0275_ VGND VGND VPWR VPWR 
+ net354
+ sky130_fd_sc_hd__dfxtp_1
X_9026_ clknet_3_4_0_wb_clk_i _0276_ VGND VGND VPWR VPWR 
+ net355
+ sky130_fd_sc_hd__dfxtp_1
X_9027_ clknet_3_4_0_wb_clk_i _0277_ VGND VGND VPWR VPWR 
+ net356
+ sky130_fd_sc_hd__dfxtp_1
X_9028_ clknet_3_5_0_wb_clk_i _0278_ VGND VGND VPWR VPWR 
+ net334
+ sky130_fd_sc_hd__dfxtp_1
X_9029_ clknet_3_5_0_wb_clk_i _0279_ VGND VGND VPWR VPWR 
+ net335
+ sky130_fd_sc_hd__dfxtp_1
X_9030_ clknet_3_5_0_wb_clk_i _0280_ VGND VGND VPWR VPWR 
+ net336
+ sky130_fd_sc_hd__dfxtp_1
X_9031_ clknet_3_5_0_wb_clk_i _0281_ VGND VGND VPWR VPWR 
+ net337
+ sky130_fd_sc_hd__dfxtp_1
X_9032_ clknet_3_5_0_wb_clk_i _0282_ VGND VGND VPWR VPWR 
+ net339
+ sky130_fd_sc_hd__dfxtp_1
X_9033_ clknet_3_7_0_wb_clk_i _0283_ VGND VGND VPWR VPWR 
+ net340
+ sky130_fd_sc_hd__dfxtp_1
X_9034_ clknet_3_7_0_wb_clk_i _0284_ VGND VGND VPWR VPWR 
+ net341
+ sky130_fd_sc_hd__dfxtp_1
X_9035_ clknet_3_5_0_wb_clk_i _0285_ VGND VGND VPWR VPWR 
+ net342
+ sky130_fd_sc_hd__dfxtp_1
X_9036_ clknet_3_7_0_wb_clk_i _0286_ VGND VGND VPWR VPWR 
+ net343
+ sky130_fd_sc_hd__dfxtp_1
X_9037_ clknet_3_7_0_wb_clk_i _0287_ VGND VGND VPWR VPWR 
+ net344
+ sky130_fd_sc_hd__dfxtp_1
X_9038_ clknet_3_7_0_wb_clk_i _0288_ VGND VGND VPWR VPWR 
+ net345
+ sky130_fd_sc_hd__dfxtp_1
X_9039_ clknet_3_5_0_wb_clk_i _0289_ VGND VGND VPWR VPWR 
+ net346
+ sky130_fd_sc_hd__dfxtp_1
X_9040_ clknet_3_7_0_wb_clk_i _0290_ VGND VGND VPWR VPWR 
+ net347
+ sky130_fd_sc_hd__dfxtp_1
X_9041_ clknet_3_7_0_wb_clk_i _0291_ VGND VGND VPWR VPWR 
+ net348
+ sky130_fd_sc_hd__dfxtp_1
X_9042_ clknet_3_7_0_wb_clk_i _0292_ VGND VGND VPWR VPWR 
+ net350
+ sky130_fd_sc_hd__dfxtp_1
X_9043_ clknet_3_7_0_wb_clk_i _0293_ VGND VGND VPWR VPWR 
+ net351
+ sky130_fd_sc_hd__dfxtp_1
X_9044_ clknet_leaf_35_csclk _0294_ VGND VGND VPWR VPWR 
+ net300
+ sky130_fd_sc_hd__dfxtp_1
X_9045_ clknet_leaf_35_csclk _0295_ VGND VGND VPWR VPWR 
+ net301
+ sky130_fd_sc_hd__dfxtp_1
X_9046_ clknet_leaf_35_csclk _0296_ VGND VGND VPWR VPWR 
+ net302
+ sky130_fd_sc_hd__dfxtp_1
X_9047_ clknet_leaf_35_csclk _0297_ VGND VGND VPWR VPWR 
+ net303
+ sky130_fd_sc_hd__dfxtp_1
X_9048_ clknet_2_1_0_mgmt_gpio_in[4] _0028_ _0216_ VGND VGND VPWR 
+ VPWR
+ \hkspi.state[0]\ sky130_fd_sc_hd__dfstp_4
X_9049_ clknet_2_1_0_mgmt_gpio_in[4] _0029_ _0217_ VGND VGND VPWR 
+ VPWR
+ \hkspi.state[1]\ sky130_fd_sc_hd__dfrtp_1
X_9050_ clknet_2_0_0_mgmt_gpio_in[4] _0030_ _0218_ VGND VGND VPWR 
+ VPWR
+ \hkspi.state[2]\ sky130_fd_sc_hd__dfrtp_2
X_9051_ clknet_2_0_0_mgmt_gpio_in[4] _0031_ _0219_ VGND VGND VPWR 
+ VPWR
+ \hkspi.state[3]\ sky130_fd_sc_hd__dfrtp_4
X_9052_ clknet_2_1_0_mgmt_gpio_in[4] _0032_ _0220_ VGND VGND VPWR 
+ VPWR
+ \hkspi.state[4]\ sky130_fd_sc_hd__dfrtp_1
X_9053_ clknet_3_3_0_wb_clk_i _0038_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_state[0]\ sky130_fd_sc_hd__dfstp_1
X_9054_ clknet_3_3_0_wb_clk_i _0039_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_state[1]\ sky130_fd_sc_hd__dfrtp_4
X_9055_ clknet_3_0_0_wb_clk_i _0040_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_state[2]\ sky130_fd_sc_hd__dfrtp_4
X_9056_ clknet_3_0_0_wb_clk_i _0041_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_state[3]\ sky130_fd_sc_hd__dfrtp_4
X_9057_ clknet_3_2_0_wb_clk_i net378 net377 VGND VGND VPWR 
+ VPWR
+ serial_resetn_pre sky130_fd_sc_hd__dfrtp_1
X_9058_ net379 _0046_ _0221_ VGND VGND VPWR 
+ VPWR
+ \hkspi.sdoenb\ sky130_fd_sc_hd__dfstp_1
X_9059_ clknet_3_6_0_wb_clk_i _0033_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[0]\ sky130_fd_sc_hd__dfstp_1
X_9060_ clknet_3_6_0_wb_clk_i _0024_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[1]\ sky130_fd_sc_hd__dfrtp_1
X_9061_ clknet_3_6_0_wb_clk_i _0025_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[2]\ sky130_fd_sc_hd__dfrtp_1
X_9062_ clknet_3_6_0_wb_clk_i _0026_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[3]\ sky130_fd_sc_hd__dfrtp_1
X_9063_ clknet_3_6_0_wb_clk_i _0027_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[4]\ sky130_fd_sc_hd__dfrtp_1
X_9064_ clknet_3_6_0_wb_clk_i _0034_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[5]\ sky130_fd_sc_hd__dfrtp_1
X_9065_ clknet_3_7_0_wb_clk_i \wbbd_state[1]\ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[6]\ sky130_fd_sc_hd__dfrtp_1
X_9066_ clknet_3_6_0_wb_clk_i _0035_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[7]\ sky130_fd_sc_hd__dfrtp_4
X_9067_ clknet_3_6_0_wb_clk_i _0036_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[8]\ sky130_fd_sc_hd__dfrtp_4
X_9068_ clknet_3_6_0_wb_clk_i _0037_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_state[9]\ sky130_fd_sc_hd__dfrtp_4
X_9069_ clknet_leaf_35_csclk _0298_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_load sky130_fd_sc_hd__dfrtp_4
X_9070_ clknet_leaf_9_csclk _0299_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][0]\ sky130_fd_sc_hd__dfstp_1
X_9071_ clknet_leaf_8_csclk _0300_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][1]\ sky130_fd_sc_hd__dfstp_1
X_9072_ clknet_leaf_8_csclk _0301_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][2]\ sky130_fd_sc_hd__dfrtp_1
X_9073_ clknet_leaf_9_csclk _0302_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][3]\ sky130_fd_sc_hd__dfrtp_2
X_9074_ clknet_leaf_9_csclk _0303_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][4]\ sky130_fd_sc_hd__dfrtp_1
X_9075_ clknet_leaf_8_csclk _0304_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][5]\ sky130_fd_sc_hd__dfrtp_1
X_9076_ clknet_leaf_9_csclk _0305_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][6]\ sky130_fd_sc_hd__dfrtp_1
X_9077_ clknet_leaf_9_csclk _0306_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][7]\ sky130_fd_sc_hd__dfrtp_1
X_9078_ clknet_leaf_35_csclk _0307_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_resetn sky130_fd_sc_hd__dfrtp_1
X_9079_ clknet_leaf_35_csclk _0308_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_data_1 sky130_fd_sc_hd__dfrtp_1
X_9080_ clknet_2_1_0_mgmt_gpio_in[4] _0309_ _0223_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pass_thru_user_delay\ sky130_fd_sc_hd__dfrtp_4
X_9081_ clknet_leaf_24_csclk _0310_ net369 VGND VGND VPWR 
+ VPWR
+ trap_output_dest sky130_fd_sc_hd__dfrtp_2
X_9082_ clknet_2_1_0_mgmt_gpio_in[4] _0311_ _0224_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[0]\ sky130_fd_sc_hd__dfrtp_2
X_9083_ clknet_2_1_0_mgmt_gpio_in[4] _0312_ _0225_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[1]\ sky130_fd_sc_hd__dfrtp_2
X_9084_ clknet_2_0_0_mgmt_gpio_in[4] _0313_ _0226_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[2]\ sky130_fd_sc_hd__dfrtp_2
X_9085_ clknet_2_2_0_mgmt_gpio_in[4] _0314_ _0227_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[3]\ sky130_fd_sc_hd__dfrtp_1
X_9086_ clknet_2_2_0_mgmt_gpio_in[4] _0315_ _0228_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[4]\ sky130_fd_sc_hd__dfrtp_2
X_9087_ clknet_2_2_0_mgmt_gpio_in[4] _0316_ _0229_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[5]\ sky130_fd_sc_hd__dfrtp_2
X_9088_ clknet_2_2_0_mgmt_gpio_in[4] _0317_ _0230_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[6]\ sky130_fd_sc_hd__dfrtp_2
X_9089_ clknet_2_2_0_mgmt_gpio_in[4] _0318_ _0231_ VGND VGND VPWR 
+ VPWR
+ \hkspi.addr[7]\ sky130_fd_sc_hd__dfrtp_1
X_9090_ clknet_2_1_0_mgmt_gpio_in[4] _0319_ _0232_ VGND VGND VPWR 
+ VPWR
+ \hkspi.count[0]\ sky130_fd_sc_hd__dfrtp_2
X_9091_ clknet_2_0_0_mgmt_gpio_in[4] _0320_ _0233_ VGND VGND VPWR 
+ VPWR
+ \hkspi.count[1]\ sky130_fd_sc_hd__dfrtp_4
X_9092_ clknet_2_0_0_mgmt_gpio_in[4] _0321_ _0234_ VGND VGND VPWR 
+ VPWR
+ \hkspi.count[2]\ sky130_fd_sc_hd__dfrtp_4
X_9093_ clknet_leaf_15_csclk _0322_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][0]\ sky130_fd_sc_hd__dfstp_1
X_9094_ clknet_leaf_15_csclk _0323_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][1]\ sky130_fd_sc_hd__dfstp_1
X_9095_ clknet_leaf_17_csclk _0324_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][2]\ sky130_fd_sc_hd__dfrtp_1
X_9096_ clknet_leaf_15_csclk _0325_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][3]\ sky130_fd_sc_hd__dfrtp_4
X_9097_ clknet_leaf_15_csclk _0326_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][4]\ sky130_fd_sc_hd__dfrtp_1
X_9098_ clknet_leaf_16_csclk _0327_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][5]\ sky130_fd_sc_hd__dfrtp_1
X_9099_ clknet_leaf_16_csclk _0328_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][6]\ sky130_fd_sc_hd__dfrtp_1
X_9100_ clknet_leaf_25_csclk _0329_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][7]\ sky130_fd_sc_hd__dfrtp_1
X_9101_ clknet_leaf_45_csclk _0330_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][8]\ sky130_fd_sc_hd__dfrtp_1
X_9102_ clknet_leaf_46_csclk _0331_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][9]\ sky130_fd_sc_hd__dfrtp_1
X_9103_ clknet_leaf_45_csclk _0332_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][10]\ sky130_fd_sc_hd__dfstp_1
X_9104_ clknet_leaf_46_csclk _0333_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][11]\ sky130_fd_sc_hd__dfrtp_1
X_9105_ clknet_leaf_45_csclk _0334_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][12]\ sky130_fd_sc_hd__dfrtp_1
X_9106_ clknet_leaf_31_csclk _0335_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][0]\ sky130_fd_sc_hd__dfstp_1
X_9107_ clknet_leaf_28_csclk _0336_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][1]\ sky130_fd_sc_hd__dfstp_1
X_9108_ clknet_leaf_31_csclk _0337_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][2]\ sky130_fd_sc_hd__dfrtp_1
X_9109_ clknet_leaf_31_csclk _0338_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][3]\ sky130_fd_sc_hd__dfrtp_1
X_9110_ clknet_leaf_32_csclk _0339_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][4]\ sky130_fd_sc_hd__dfrtp_1
X_9111_ clknet_leaf_31_csclk _0340_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][5]\ sky130_fd_sc_hd__dfrtp_1
X_9112_ clknet_leaf_31_csclk _0341_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][6]\ sky130_fd_sc_hd__dfrtp_1
X_9113_ clknet_leaf_28_csclk _0342_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[4][7]\ sky130_fd_sc_hd__dfrtp_1
X_9114_ clknet_leaf_41_csclk _0343_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][8]\ sky130_fd_sc_hd__dfrtp_1
X_9115_ clknet_leaf_30_csclk _0344_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][9]\ sky130_fd_sc_hd__dfrtp_1
X_9116_ clknet_leaf_41_csclk _0345_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][10]\ sky130_fd_sc_hd__dfstp_1
X_9117_ clknet_leaf_40_csclk _0346_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][11]\ sky130_fd_sc_hd__dfrtp_1
X_9118_ clknet_leaf_41_csclk _0347_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][12]\ sky130_fd_sc_hd__dfrtp_1
X_9119_ clknet_3_6_0_wb_clk_i _0348_ net196 VGND VGND VPWR 
+ VPWR
+ net326 sky130_fd_sc_hd__dfrtp_4
X_9120_ clknet_leaf_39_csclk _0349_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][8]\ sky130_fd_sc_hd__dfrtp_1
X_9121_ clknet_leaf_39_csclk _0350_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][9]\ sky130_fd_sc_hd__dfrtp_1
X_9122_ clknet_leaf_40_csclk _0351_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][10]\ sky130_fd_sc_hd__dfstp_1
X_9123_ clknet_leaf_39_csclk _0352_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][11]\ sky130_fd_sc_hd__dfrtp_1
X_9124_ clknet_leaf_39_csclk _0353_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][12]\ sky130_fd_sc_hd__dfrtp_1
X_9125_ clknet_leaf_31_csclk _0354_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][0]\ sky130_fd_sc_hd__dfstp_1
X_9126_ clknet_leaf_30_csclk _0355_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][1]\ sky130_fd_sc_hd__dfstp_1
X_9127_ clknet_leaf_31_csclk _0356_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][2]\ sky130_fd_sc_hd__dfrtp_1
X_9128_ clknet_leaf_31_csclk _0357_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][3]\ sky130_fd_sc_hd__dfrtp_1
X_9129_ clknet_leaf_30_csclk _0358_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][4]\ sky130_fd_sc_hd__dfrtp_1
X_9130_ clknet_leaf_31_csclk _0359_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][5]\ sky130_fd_sc_hd__dfrtp_1
X_9131_ clknet_leaf_31_csclk _0360_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][6]\ sky130_fd_sc_hd__dfrtp_1
X_9132_ clknet_leaf_31_csclk _0361_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[6][7]\ sky130_fd_sc_hd__dfrtp_1
X_9133_ clknet_leaf_7_csclk _0362_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][8]\ sky130_fd_sc_hd__dfrtp_1
X_9134_ clknet_leaf_8_csclk _0363_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][9]\ sky130_fd_sc_hd__dfrtp_1
X_9135_ clknet_leaf_7_csclk _0364_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][10]\ sky130_fd_sc_hd__dfstp_1
X_9136_ clknet_leaf_7_csclk _0365_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][11]\ sky130_fd_sc_hd__dfrtp_1
X_9137_ clknet_leaf_7_csclk _0366_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][12]\ sky130_fd_sc_hd__dfrtp_1
X_9138_ clknet_3_0_0_wb_clk_i _0367_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[0]\ sky130_fd_sc_hd__dfrtp_1
X_9139_ clknet_3_3_0_wb_clk_i _0368_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[1]\ sky130_fd_sc_hd__dfrtp_1
X_9140_ clknet_3_3_0_wb_clk_i _0369_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[2]\ sky130_fd_sc_hd__dfrtp_1
X_9141_ clknet_3_3_0_wb_clk_i _0370_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[3]\ sky130_fd_sc_hd__dfrtp_1
X_9142_ clknet_3_3_0_wb_clk_i _0371_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[4]\ sky130_fd_sc_hd__dfrtp_1
X_9143_ clknet_3_0_0_wb_clk_i _0372_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[5]\ sky130_fd_sc_hd__dfrtp_1
X_9144_ clknet_3_3_0_wb_clk_i _0373_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[6]\ sky130_fd_sc_hd__dfrtp_1
X_9145_ clknet_3_0_0_wb_clk_i _0374_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[7]\ sky130_fd_sc_hd__dfrtp_1
X_9146_ clknet_3_2_0_wb_clk_i _0375_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[8]\ sky130_fd_sc_hd__dfrtp_1
X_9147_ clknet_3_2_0_wb_clk_i _0376_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[9]\ sky130_fd_sc_hd__dfrtp_1
X_9148_ clknet_3_2_0_wb_clk_i _0377_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[10]\ sky130_fd_sc_hd__dfrtp_1
X_9149_ clknet_3_2_0_wb_clk_i _0378_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[11]\ sky130_fd_sc_hd__dfrtp_1
X_9150_ clknet_3_2_0_wb_clk_i _0379_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_2[12]\ sky130_fd_sc_hd__dfrtp_1
X_9151_ clknet_leaf_28_csclk _0380_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][0]\ sky130_fd_sc_hd__dfstp_1
X_9152_ clknet_leaf_27_csclk _0381_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][1]\ sky130_fd_sc_hd__dfstp_1
X_9153_ clknet_leaf_27_csclk _0382_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][2]\ sky130_fd_sc_hd__dfrtp_1
X_9154_ clknet_leaf_32_csclk _0383_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][3]\ sky130_fd_sc_hd__dfrtp_1
X_9155_ clknet_leaf_32_csclk _0384_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][4]\ sky130_fd_sc_hd__dfrtp_1
X_9156_ clknet_leaf_32_csclk _0385_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][5]\ sky130_fd_sc_hd__dfrtp_1
X_9157_ clknet_leaf_28_csclk _0386_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][6]\ sky130_fd_sc_hd__dfrtp_1
X_9158_ clknet_leaf_32_csclk _0387_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[7][7]\ sky130_fd_sc_hd__dfrtp_1
X_9159_ clknet_leaf_8_csclk _0388_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][8]\ sky130_fd_sc_hd__dfrtp_1
X_9160_ clknet_leaf_8_csclk _0389_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][9]\ sky130_fd_sc_hd__dfrtp_1
X_9161_ clknet_leaf_13_csclk _0390_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][10]\ sky130_fd_sc_hd__dfstp_1
X_9162_ clknet_leaf_8_csclk _0391_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][11]\ sky130_fd_sc_hd__dfrtp_1
X_9163_ clknet_leaf_13_csclk _0392_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][12]\ sky130_fd_sc_hd__dfrtp_1
X_9164_ clknet_3_0_0_wb_clk_i _0393_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[0]\ sky130_fd_sc_hd__dfrtp_1
X_9165_ clknet_3_0_0_wb_clk_i _0394_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[1]\ sky130_fd_sc_hd__dfrtp_1
X_9166_ clknet_3_0_0_wb_clk_i _0395_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[2]\ sky130_fd_sc_hd__dfrtp_1
X_9167_ clknet_3_0_0_wb_clk_i _0396_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[3]\ sky130_fd_sc_hd__dfrtp_1
X_9168_ clknet_3_0_0_wb_clk_i _0397_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[4]\ sky130_fd_sc_hd__dfrtp_1
X_9169_ clknet_3_0_0_wb_clk_i _0398_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[5]\ sky130_fd_sc_hd__dfrtp_1
X_9170_ clknet_3_0_0_wb_clk_i _0399_ net376 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[6]\ sky130_fd_sc_hd__dfrtp_1
X_9171_ clknet_3_2_0_wb_clk_i _0400_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[7]\ sky130_fd_sc_hd__dfrtp_1
X_9172_ clknet_3_0_0_wb_clk_i _0401_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[8]\ sky130_fd_sc_hd__dfrtp_1
X_9173_ clknet_3_2_0_wb_clk_i _0402_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[9]\ sky130_fd_sc_hd__dfrtp_1
X_9174_ clknet_3_2_0_wb_clk_i _0403_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[10]\ sky130_fd_sc_hd__dfrtp_1
X_9175_ clknet_3_2_0_wb_clk_i _0404_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[11]\ sky130_fd_sc_hd__dfrtp_1
X_9176_ clknet_3_2_0_wb_clk_i _0405_ net377 VGND VGND VPWR 
+ VPWR
+ \serial_data_staging_1[12]\ sky130_fd_sc_hd__dfrtp_1
X_9177_ clknet_leaf_26_csclk _0406_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][0]\ sky130_fd_sc_hd__dfstp_1
X_9178_ clknet_leaf_26_csclk _0407_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][1]\ sky130_fd_sc_hd__dfstp_1
X_9179_ clknet_leaf_25_csclk _0408_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][2]\ sky130_fd_sc_hd__dfrtp_1
X_9180_ clknet_leaf_26_csclk _0409_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][3]\ sky130_fd_sc_hd__dfrtp_4
X_9181_ clknet_leaf_26_csclk _0410_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][4]\ sky130_fd_sc_hd__dfrtp_1
X_9182_ clknet_leaf_25_csclk _0411_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][5]\ sky130_fd_sc_hd__dfrtp_1
X_9183_ clknet_leaf_26_csclk _0412_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][6]\ sky130_fd_sc_hd__dfrtp_1
X_9184_ clknet_leaf_26_csclk _0413_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[8][7]\ sky130_fd_sc_hd__dfrtp_1
X_9185_ clknet_leaf_39_csclk _0414_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][8]\ sky130_fd_sc_hd__dfrtp_1
X_9186_ clknet_leaf_43_csclk _0415_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][9]\ sky130_fd_sc_hd__dfrtp_1
X_9187_ clknet_leaf_38_csclk _0416_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][10]\ sky130_fd_sc_hd__dfstp_1
X_9188_ clknet_leaf_43_csclk _0417_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][11]\ sky130_fd_sc_hd__dfrtp_1
X_9189_ clknet_leaf_39_csclk _0418_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][12]\ sky130_fd_sc_hd__dfrtp_1
X_9190_ clknet_leaf_27_csclk _0419_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][0]\ sky130_fd_sc_hd__dfstp_1
X_9191_ clknet_leaf_28_csclk _0420_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][1]\ sky130_fd_sc_hd__dfstp_1
X_9192_ clknet_leaf_28_csclk _0421_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][2]\ sky130_fd_sc_hd__dfrtp_1
X_9193_ clknet_leaf_28_csclk _0422_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][3]\ sky130_fd_sc_hd__dfrtp_1
X_9194_ clknet_leaf_28_csclk _0423_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][4]\ sky130_fd_sc_hd__dfrtp_1
X_9195_ clknet_leaf_29_csclk _0424_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][5]\ sky130_fd_sc_hd__dfrtp_1
X_9196_ clknet_leaf_29_csclk _0425_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][6]\ sky130_fd_sc_hd__dfrtp_1
X_9197_ clknet_leaf_29_csclk _0426_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[9][7]\ sky130_fd_sc_hd__dfrtp_1
X_9198_ clknet_leaf_6_csclk _0427_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][8]\ sky130_fd_sc_hd__dfrtp_1
X_9199_ clknet_leaf_5_csclk _0428_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][9]\ sky130_fd_sc_hd__dfrtp_1
X_9200_ clknet_leaf_5_csclk _0429_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][10]\ sky130_fd_sc_hd__dfstp_1
X_9201_ clknet_leaf_5_csclk _0430_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][11]\ sky130_fd_sc_hd__dfrtp_1
X_9202_ clknet_leaf_6_csclk _0431_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][12]\ sky130_fd_sc_hd__dfrtp_1
X_9203_ clknet_3_0_0_wb_clk_i _0432_ net376 VGND VGND VPWR 
+ VPWR
+ serial_busy sky130_fd_sc_hd__dfrtp_1
X_9204_ clknet_leaf_25_csclk _0433_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][0]\ sky130_fd_sc_hd__dfstp_1
X_9205_ clknet_leaf_26_csclk _0434_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][1]\ sky130_fd_sc_hd__dfstp_1
X_9206_ clknet_leaf_25_csclk _0435_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][2]\ sky130_fd_sc_hd__dfrtp_1
X_9207_ clknet_leaf_24_csclk _0436_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][3]\ sky130_fd_sc_hd__dfrtp_2
X_9208_ clknet_leaf_24_csclk _0437_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][4]\ sky130_fd_sc_hd__dfrtp_1
X_9209_ clknet_leaf_25_csclk _0438_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][5]\ sky130_fd_sc_hd__dfrtp_1
X_9210_ clknet_leaf_25_csclk _0439_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][6]\ sky130_fd_sc_hd__dfrtp_1
X_9211_ clknet_leaf_26_csclk _0440_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[10][7]\ sky130_fd_sc_hd__dfrtp_1
X_9212_ clknet_leaf_39_csclk _0441_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][8]\ sky130_fd_sc_hd__dfrtp_1
X_9213_ clknet_leaf_43_csclk _0442_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][9]\ sky130_fd_sc_hd__dfrtp_1
X_9214_ clknet_leaf_39_csclk _0443_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][10]\ sky130_fd_sc_hd__dfstp_1
X_9215_ clknet_leaf_43_csclk _0444_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][11]\ sky130_fd_sc_hd__dfrtp_1
X_9216_ clknet_leaf_39_csclk _0445_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][12]\ sky130_fd_sc_hd__dfrtp_1
X_9217_ clknet_3_2_0_wb_clk_i _0446_ net377 VGND VGND VPWR 
+ VPWR
+ serial_load_pre sky130_fd_sc_hd__dfrtp_1
X_9218_ clknet_leaf_31_csclk _0447_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][0]\ sky130_fd_sc_hd__dfstp_1
X_9219_ clknet_leaf_32_csclk _0448_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][1]\ sky130_fd_sc_hd__dfstp_1
X_9220_ clknet_leaf_32_csclk _0449_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][2]\ sky130_fd_sc_hd__dfrtp_1
X_9221_ clknet_leaf_32_csclk _0450_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][3]\ sky130_fd_sc_hd__dfrtp_1
X_9222_ clknet_leaf_32_csclk _0451_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][4]\ sky130_fd_sc_hd__dfrtp_1
X_9223_ clknet_leaf_32_csclk _0452_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][5]\ sky130_fd_sc_hd__dfrtp_1
X_9224_ clknet_leaf_32_csclk _0453_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][6]\ sky130_fd_sc_hd__dfrtp_1
X_9225_ clknet_leaf_32_csclk _0454_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[11][7]\ sky130_fd_sc_hd__dfrtp_1
X_9226_ clknet_leaf_6_csclk _0455_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][8]\ sky130_fd_sc_hd__dfrtp_1
X_9227_ clknet_leaf_6_csclk _0456_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][9]\ sky130_fd_sc_hd__dfrtp_1
X_9228_ clknet_leaf_6_csclk _0457_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][10]\ sky130_fd_sc_hd__dfstp_1
X_9229_ clknet_leaf_6_csclk _0458_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][11]\ sky130_fd_sc_hd__dfrtp_1
X_9230_ clknet_leaf_6_csclk _0459_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][12]\ sky130_fd_sc_hd__dfrtp_1
X_9231_ clknet_leaf_17_csclk _0460_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][0]\ sky130_fd_sc_hd__dfstp_1
X_9232_ clknet_leaf_17_csclk _0461_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][1]\ sky130_fd_sc_hd__dfstp_1
X_9233_ clknet_leaf_17_csclk _0462_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][2]\ sky130_fd_sc_hd__dfrtp_1
X_9234_ clknet_leaf_21_csclk _0463_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][3]\ sky130_fd_sc_hd__dfrtp_2
X_9235_ clknet_leaf_17_csclk _0464_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][4]\ sky130_fd_sc_hd__dfrtp_1
X_9236_ clknet_leaf_21_csclk _0465_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][5]\ sky130_fd_sc_hd__dfrtp_1
X_9237_ clknet_leaf_20_csclk _0466_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][6]\ sky130_fd_sc_hd__dfrtp_1
X_9238_ clknet_leaf_21_csclk _0467_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[12][7]\ sky130_fd_sc_hd__dfrtp_1
X_9239_ clknet_3_3_0_wb_clk_i _0468_ net377 VGND VGND VPWR 
+ VPWR
+ serial_clock_pre sky130_fd_sc_hd__dfrtp_2
X_9240_ clknet_leaf_5_csclk _0469_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][8]\ sky130_fd_sc_hd__dfrtp_1
X_9241_ clknet_leaf_5_csclk _0470_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][9]\ sky130_fd_sc_hd__dfrtp_1
X_9242_ clknet_leaf_5_csclk _0471_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][10]\ sky130_fd_sc_hd__dfstp_1
X_9243_ clknet_leaf_5_csclk _0472_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][11]\ sky130_fd_sc_hd__dfrtp_1
X_9244_ clknet_leaf_5_csclk _0473_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][12]\ sky130_fd_sc_hd__dfrtp_1
X_9245_ clknet_3_3_0_wb_clk_i _0474_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[0]\ sky130_fd_sc_hd__dfstp_2
X_9246_ clknet_3_3_0_wb_clk_i _0475_ net370 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[1]\ sky130_fd_sc_hd__dfstp_2
X_9247_ clknet_3_3_0_wb_clk_i _0476_ net370 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[2]\ sky130_fd_sc_hd__dfrtp_1
X_9248_ clknet_3_3_0_wb_clk_i _0477_ net370 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[3]\ sky130_fd_sc_hd__dfrtp_2
X_9249_ clknet_3_3_0_wb_clk_i _0478_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[4]\ sky130_fd_sc_hd__dfstp_1
X_9250_ clknet_3_3_0_wb_clk_i _0479_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_2[5]\ sky130_fd_sc_hd__dfrtp_1
X_9251_ clknet_3_3_0_wb_clk_i _0480_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_1[0]\ sky130_fd_sc_hd__dfrtp_4
X_9252_ clknet_3_3_0_wb_clk_i _0481_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_1[1]\ sky130_fd_sc_hd__dfstp_1
X_9253_ clknet_3_1_0_wb_clk_i _0482_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_1[2]\ sky130_fd_sc_hd__dfrtp_2
X_9254_ clknet_3_1_0_wb_clk_i _0483_ net376 VGND VGND VPWR 
+ VPWR
+ \pad_count_1[3]\ sky130_fd_sc_hd__dfrtp_1
X_9255_ clknet_3_3_0_wb_clk_i _0484_ net370 VGND VGND VPWR 
+ VPWR
+ \pad_count_1[4]\ sky130_fd_sc_hd__dfstp_4
X_9256_ clknet_leaf_22_csclk _0485_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][0]\ sky130_fd_sc_hd__dfstp_1
X_9257_ clknet_leaf_22_csclk _0486_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][1]\ sky130_fd_sc_hd__dfstp_1
X_9258_ clknet_leaf_22_csclk _0487_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][2]\ sky130_fd_sc_hd__dfrtp_1
X_9259_ clknet_leaf_22_csclk _0488_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][3]\ sky130_fd_sc_hd__dfrtp_2
X_9260_ clknet_leaf_22_csclk _0489_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][4]\ sky130_fd_sc_hd__dfrtp_1
X_9261_ clknet_leaf_22_csclk _0490_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][5]\ sky130_fd_sc_hd__dfrtp_1
X_9262_ clknet_leaf_22_csclk _0491_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][6]\ sky130_fd_sc_hd__dfrtp_1
X_9263_ clknet_leaf_22_csclk _0492_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[13][7]\ sky130_fd_sc_hd__dfrtp_1
X_9264_ clknet_leaf_7_csclk _0493_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][8]\ sky130_fd_sc_hd__dfrtp_1
X_9265_ clknet_leaf_5_csclk _0494_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][9]\ sky130_fd_sc_hd__dfrtp_1
X_9266_ clknet_leaf_7_csclk _0495_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][10]\ sky130_fd_sc_hd__dfstp_1
X_9267_ clknet_leaf_7_csclk _0496_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][11]\ sky130_fd_sc_hd__dfrtp_1
X_9268_ clknet_leaf_7_csclk _0497_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][12]\ sky130_fd_sc_hd__dfrtp_1
X_9269_ clknet_leaf_12_csclk _0498_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][0]\ sky130_fd_sc_hd__dfstp_1
X_9270_ clknet_leaf_12_csclk _0499_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][1]\ sky130_fd_sc_hd__dfstp_1
X_9271_ clknet_leaf_12_csclk _0500_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][2]\ sky130_fd_sc_hd__dfrtp_1
X_9272_ clknet_leaf_16_csclk _0501_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][3]\ sky130_fd_sc_hd__dfrtp_1
X_9273_ clknet_leaf_12_csclk _0502_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][4]\ sky130_fd_sc_hd__dfrtp_1
X_9274_ clknet_leaf_21_csclk _0503_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][5]\ sky130_fd_sc_hd__dfrtp_1
X_9275_ clknet_leaf_21_csclk _0504_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][6]\ sky130_fd_sc_hd__dfrtp_1
X_9276_ clknet_leaf_20_csclk _0505_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[14][7]\ sky130_fd_sc_hd__dfrtp_1
X_9277_ clknet_3_3_0_wb_clk_i _0506_ net377 VGND VGND VPWR 
+ VPWR
+ \xfer_count[0]\ sky130_fd_sc_hd__dfrtp_2
X_9278_ clknet_3_3_0_wb_clk_i _0507_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_count[1]\ sky130_fd_sc_hd__dfrtp_1
X_9279_ clknet_3_2_0_wb_clk_i _0508_ net376 VGND VGND VPWR 
+ VPWR
+ \xfer_count[2]\ sky130_fd_sc_hd__dfrtp_1
X_9280_ clknet_3_2_0_wb_clk_i _0509_ net377 VGND VGND VPWR 
+ VPWR
+ \xfer_count[3]\ sky130_fd_sc_hd__dfrtp_1
X_9281_ clknet_leaf_9_csclk _0510_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][8]\ sky130_fd_sc_hd__dfrtp_1
X_9282_ clknet_leaf_9_csclk _0511_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][9]\ sky130_fd_sc_hd__dfrtp_1
X_9283_ clknet_leaf_9_csclk _0512_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][10]\ sky130_fd_sc_hd__dfstp_1
X_9284_ clknet_leaf_8_csclk _0513_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][11]\ sky130_fd_sc_hd__dfrtp_1
X_9285_ clknet_leaf_9_csclk _0514_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][12]\ sky130_fd_sc_hd__dfrtp_1
X_9286_ clknet_leaf_18_csclk _0515_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][0]\ sky130_fd_sc_hd__dfstp_1
X_9287_ clknet_leaf_18_csclk _0516_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][1]\ sky130_fd_sc_hd__dfstp_1
X_9288_ clknet_leaf_18_csclk _0517_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][2]\ sky130_fd_sc_hd__dfrtp_1
X_9289_ clknet_leaf_20_csclk _0518_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][3]\ sky130_fd_sc_hd__dfrtp_1
X_9290_ clknet_leaf_18_csclk _0519_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][4]\ sky130_fd_sc_hd__dfrtp_1
X_9291_ clknet_leaf_20_csclk _0520_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][5]\ sky130_fd_sc_hd__dfrtp_1
X_9292_ clknet_leaf_20_csclk _0521_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][6]\ sky130_fd_sc_hd__dfrtp_1
X_9293_ clknet_leaf_20_csclk _0522_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][7]\ sky130_fd_sc_hd__dfrtp_1
X_9294_ clknet_leaf_21_csclk _0523_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][0]\ sky130_fd_sc_hd__dfstp_1
X_9295_ clknet_leaf_21_csclk _0524_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][1]\ sky130_fd_sc_hd__dfstp_1
X_9296_ clknet_leaf_24_csclk _0525_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][2]\ sky130_fd_sc_hd__dfrtp_1
X_9297_ clknet_leaf_24_csclk _0526_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][3]\ sky130_fd_sc_hd__dfrtp_2
X_9298_ clknet_leaf_24_csclk _0527_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][4]\ sky130_fd_sc_hd__dfrtp_1
X_9299_ clknet_leaf_21_csclk _0528_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][5]\ sky130_fd_sc_hd__dfrtp_1
X_9300_ clknet_leaf_24_csclk _0529_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][6]\ sky130_fd_sc_hd__dfrtp_1
X_9301_ clknet_leaf_24_csclk _0530_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[15][7]\ sky130_fd_sc_hd__dfrtp_1
X_9302_ clknet_leaf_6_csclk _0531_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][8]\ sky130_fd_sc_hd__dfrtp_1
X_9303_ clknet_leaf_6_csclk _0532_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][9]\ sky130_fd_sc_hd__dfrtp_1
X_9304_ clknet_leaf_6_csclk _0533_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][10]\ sky130_fd_sc_hd__dfrtp_1
X_9305_ clknet_leaf_6_csclk _0534_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][11]\ sky130_fd_sc_hd__dfstp_1
X_9306_ clknet_leaf_6_csclk _0535_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[37][12]\ sky130_fd_sc_hd__dfstp_1
X_9307_ clknet_leaf_5_csclk _0536_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][8]\ sky130_fd_sc_hd__dfrtp_1
X_9308_ clknet_leaf_5_csclk _0537_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][9]\ sky130_fd_sc_hd__dfrtp_1
X_9309_ clknet_leaf_5_csclk _0538_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][10]\ sky130_fd_sc_hd__dfstp_1
X_9310_ clknet_leaf_5_csclk _0539_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][11]\ sky130_fd_sc_hd__dfrtp_1
X_9311_ clknet_leaf_5_csclk _0540_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][12]\ sky130_fd_sc_hd__dfrtp_1
X_9312_ clknet_leaf_14_csclk _0541_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][0]\ sky130_fd_sc_hd__dfstp_1
X_9313_ clknet_leaf_14_csclk _0542_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][1]\ sky130_fd_sc_hd__dfstp_1
X_9314_ clknet_leaf_14_csclk _0543_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][2]\ sky130_fd_sc_hd__dfrtp_1
X_9315_ clknet_leaf_12_csclk _0544_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][3]\ sky130_fd_sc_hd__dfrtp_1
X_9316_ clknet_leaf_14_csclk _0545_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][4]\ sky130_fd_sc_hd__dfrtp_1
X_9317_ clknet_leaf_15_csclk _0546_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][5]\ sky130_fd_sc_hd__dfrtp_1
X_9318_ clknet_leaf_17_csclk _0547_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][6]\ sky130_fd_sc_hd__dfrtp_1
X_9319_ clknet_leaf_16_csclk _0548_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][7]\ sky130_fd_sc_hd__dfrtp_1
X_9320_ clknet_leaf_26_csclk _0549_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][0]\ sky130_fd_sc_hd__dfstp_1
X_9321_ clknet_leaf_27_csclk _0550_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][1]\ sky130_fd_sc_hd__dfstp_1
X_9322_ clknet_leaf_27_csclk _0551_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][2]\ sky130_fd_sc_hd__dfrtp_1
X_9323_ clknet_leaf_26_csclk _0552_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][3]\ sky130_fd_sc_hd__dfrtp_4
X_9324_ clknet_leaf_27_csclk _0553_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][4]\ sky130_fd_sc_hd__dfrtp_1
X_9325_ clknet_leaf_26_csclk _0554_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][5]\ sky130_fd_sc_hd__dfrtp_1
X_9326_ clknet_leaf_27_csclk _0555_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][6]\ sky130_fd_sc_hd__dfrtp_1
X_9327_ clknet_leaf_27_csclk _0556_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[16][7]\ sky130_fd_sc_hd__dfrtp_1
X_9328_ clknet_leaf_4_csclk _0557_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][8]\ sky130_fd_sc_hd__dfrtp_1
X_9329_ clknet_2_0_0_csclk _0558_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][9]\ sky130_fd_sc_hd__dfrtp_1
X_9330_ clknet_leaf_47_csclk _0559_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][10]\ sky130_fd_sc_hd__dfrtp_1
X_9331_ clknet_leaf_3_csclk _0560_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][11]\ sky130_fd_sc_hd__dfstp_1
X_9332_ clknet_leaf_0_csclk _0561_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[36][12]\ sky130_fd_sc_hd__dfstp_1
X_9333_ clknet_leaf_12_csclk _0562_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][8]\ sky130_fd_sc_hd__dfrtp_1
X_9334_ clknet_leaf_13_csclk _0563_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][9]\ sky130_fd_sc_hd__dfrtp_1
X_9335_ clknet_leaf_12_csclk _0564_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][10]\ sky130_fd_sc_hd__dfstp_1
X_9336_ clknet_leaf_13_csclk _0565_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][11]\ sky130_fd_sc_hd__dfrtp_1
X_9337_ clknet_leaf_13_csclk _0566_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][12]\ sky130_fd_sc_hd__dfrtp_1
X_9338_ clknet_leaf_12_csclk _0567_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][0]\ sky130_fd_sc_hd__dfstp_1
X_9339_ clknet_leaf_17_csclk _0568_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][1]\ sky130_fd_sc_hd__dfstp_1
X_9340_ clknet_leaf_12_csclk _0569_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][2]\ sky130_fd_sc_hd__dfrtp_1
X_9341_ clknet_leaf_16_csclk _0570_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][3]\ sky130_fd_sc_hd__dfrtp_1
X_9342_ clknet_leaf_17_csclk _0571_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][4]\ sky130_fd_sc_hd__dfrtp_1
X_9343_ clknet_leaf_16_csclk _0572_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][5]\ sky130_fd_sc_hd__dfrtp_1
X_9344_ clknet_leaf_16_csclk _0573_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][6]\ sky130_fd_sc_hd__dfrtp_1
X_9345_ clknet_leaf_21_csclk _0574_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][7]\ sky130_fd_sc_hd__dfrtp_1
X_9346_ clknet_leaf_27_csclk _0575_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][0]\ sky130_fd_sc_hd__dfstp_1
X_9347_ clknet_leaf_27_csclk _0576_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][1]\ sky130_fd_sc_hd__dfstp_1
X_9348_ clknet_leaf_27_csclk _0577_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][2]\ sky130_fd_sc_hd__dfrtp_1
X_9349_ clknet_leaf_26_csclk _0578_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][3]\ sky130_fd_sc_hd__dfrtp_4
X_9350_ clknet_leaf_27_csclk _0579_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][4]\ sky130_fd_sc_hd__dfrtp_1
X_9351_ clknet_leaf_26_csclk _0580_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][5]\ sky130_fd_sc_hd__dfrtp_1
X_9352_ clknet_leaf_27_csclk _0581_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][6]\ sky130_fd_sc_hd__dfrtp_1
X_9353_ clknet_leaf_28_csclk _0582_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[17][7]\ sky130_fd_sc_hd__dfrtp_1
X_9354_ clknet_leaf_7_csclk _0583_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][8]\ sky130_fd_sc_hd__dfrtp_1
X_9355_ clknet_leaf_8_csclk _0584_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][9]\ sky130_fd_sc_hd__dfrtp_1
X_9356_ clknet_leaf_8_csclk _0585_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][10]\ sky130_fd_sc_hd__dfstp_1
X_9357_ clknet_leaf_8_csclk _0586_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][11]\ sky130_fd_sc_hd__dfrtp_1
X_9358_ clknet_leaf_8_csclk _0587_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[35][12]\ sky130_fd_sc_hd__dfrtp_1
X_9359_ clknet_leaf_1_csclk _0588_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][8]\ sky130_fd_sc_hd__dfrtp_1
X_9360_ clknet_leaf_3_csclk _0589_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][9]\ sky130_fd_sc_hd__dfrtp_1
X_9361_ clknet_leaf_0_csclk _0590_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][10]\ sky130_fd_sc_hd__dfstp_1
X_9362_ clknet_leaf_2_csclk _0591_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][11]\ sky130_fd_sc_hd__dfrtp_1
X_9363_ clknet_leaf_3_csclk _0592_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][12]\ sky130_fd_sc_hd__dfrtp_1
X_9364_ clknet_leaf_17_csclk _0593_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][0]\ sky130_fd_sc_hd__dfstp_1
X_9365_ clknet_leaf_17_csclk _0594_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][1]\ sky130_fd_sc_hd__dfstp_1
X_9366_ clknet_leaf_17_csclk _0595_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][2]\ sky130_fd_sc_hd__dfrtp_1
X_9367_ clknet_leaf_21_csclk _0596_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][3]\ sky130_fd_sc_hd__dfrtp_1
X_9368_ clknet_leaf_17_csclk _0597_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][4]\ sky130_fd_sc_hd__dfrtp_1
X_9369_ clknet_leaf_21_csclk _0598_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][5]\ sky130_fd_sc_hd__dfrtp_1
X_9370_ clknet_leaf_21_csclk _0599_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][6]\ sky130_fd_sc_hd__dfrtp_1
X_9371_ clknet_leaf_21_csclk _0600_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][7]\ sky130_fd_sc_hd__dfrtp_1
X_9372_ clknet_leaf_31_csclk _0601_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][0]\ sky130_fd_sc_hd__dfstp_1
X_9373_ clknet_leaf_31_csclk _0602_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][1]\ sky130_fd_sc_hd__dfstp_1
X_9374_ clknet_leaf_31_csclk _0603_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][2]\ sky130_fd_sc_hd__dfrtp_1
X_9375_ clknet_leaf_31_csclk _0604_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][3]\ sky130_fd_sc_hd__dfrtp_4
X_9376_ clknet_leaf_31_csclk _0605_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][4]\ sky130_fd_sc_hd__dfrtp_1
X_9377_ clknet_leaf_28_csclk _0606_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][5]\ sky130_fd_sc_hd__dfrtp_1
X_9378_ clknet_leaf_28_csclk _0607_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][6]\ sky130_fd_sc_hd__dfrtp_1
X_9379_ clknet_leaf_31_csclk _0608_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[18][7]\ sky130_fd_sc_hd__dfrtp_1
X_9380_ clknet_leaf_4_csclk _0609_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][8]\ sky130_fd_sc_hd__dfrtp_1
X_9381_ clknet_leaf_3_csclk _0610_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][9]\ sky130_fd_sc_hd__dfrtp_1
X_9382_ clknet_leaf_3_csclk _0611_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][10]\ sky130_fd_sc_hd__dfstp_1
X_9383_ clknet_leaf_3_csclk _0612_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][11]\ sky130_fd_sc_hd__dfrtp_1
X_9384_ clknet_leaf_3_csclk _0613_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[34][12]\ sky130_fd_sc_hd__dfrtp_1
X_9385_ clknet_leaf_46_csclk _0614_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][8]\ sky130_fd_sc_hd__dfrtp_1
X_9386_ clknet_leaf_45_csclk _0615_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][9]\ sky130_fd_sc_hd__dfrtp_1
X_9387_ clknet_leaf_46_csclk _0616_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][10]\ sky130_fd_sc_hd__dfstp_1
X_9388_ clknet_leaf_46_csclk _0617_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][11]\ sky130_fd_sc_hd__dfrtp_1
X_9389_ clknet_leaf_46_csclk _0618_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][12]\ sky130_fd_sc_hd__dfrtp_1
X_9390_ clknet_leaf_18_csclk _0619_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][0]\ sky130_fd_sc_hd__dfstp_1
X_9391_ clknet_leaf_18_csclk _0620_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][1]\ sky130_fd_sc_hd__dfstp_1
X_9392_ clknet_leaf_18_csclk _0621_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][2]\ sky130_fd_sc_hd__dfrtp_1
X_9393_ clknet_leaf_19_csclk _0622_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][3]\ sky130_fd_sc_hd__dfrtp_1
X_9394_ clknet_leaf_18_csclk _0623_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][4]\ sky130_fd_sc_hd__dfrtp_1
X_9395_ clknet_leaf_19_csclk _0624_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][5]\ sky130_fd_sc_hd__dfrtp_1
X_9396_ clknet_leaf_19_csclk _0625_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][6]\ sky130_fd_sc_hd__dfrtp_1
X_9397_ clknet_leaf_19_csclk _0626_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][7]\ sky130_fd_sc_hd__dfrtp_1
X_9398_ clknet_leaf_43_csclk _0627_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][0]\ sky130_fd_sc_hd__dfstp_1
X_9399_ clknet_leaf_43_csclk _0628_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][1]\ sky130_fd_sc_hd__dfstp_1
X_9400_ clknet_leaf_43_csclk _0629_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][2]\ sky130_fd_sc_hd__dfrtp_1
X_9401_ clknet_leaf_43_csclk _0630_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][3]\ sky130_fd_sc_hd__dfrtp_2
X_9402_ clknet_leaf_43_csclk _0631_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][4]\ sky130_fd_sc_hd__dfrtp_1
X_9403_ clknet_leaf_43_csclk _0632_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][5]\ sky130_fd_sc_hd__dfrtp_1
X_9404_ clknet_leaf_43_csclk _0633_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][6]\ sky130_fd_sc_hd__dfrtp_4
X_9405_ clknet_leaf_43_csclk _0634_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[19][7]\ sky130_fd_sc_hd__dfrtp_1
X_9406_ clknet_leaf_1_csclk _0635_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][8]\ sky130_fd_sc_hd__dfrtp_1
X_9407_ clknet_leaf_1_csclk _0636_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][9]\ sky130_fd_sc_hd__dfrtp_1
X_9408_ clknet_leaf_1_csclk _0637_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][10]\ sky130_fd_sc_hd__dfstp_1
X_9409_ clknet_leaf_1_csclk _0638_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][11]\ sky130_fd_sc_hd__dfrtp_1
X_9410_ clknet_leaf_2_csclk _0639_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[33][12]\ sky130_fd_sc_hd__dfrtp_1
X_9411_ clknet_leaf_2_csclk _0640_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][8]\ sky130_fd_sc_hd__dfrtp_1
X_9412_ clknet_leaf_1_csclk _0641_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][9]\ sky130_fd_sc_hd__dfrtp_1
X_9413_ clknet_leaf_2_csclk _0642_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][10]\ sky130_fd_sc_hd__dfstp_1
X_9414_ clknet_leaf_2_csclk _0643_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][11]\ sky130_fd_sc_hd__dfrtp_1
X_9415_ clknet_leaf_2_csclk _0644_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][12]\ sky130_fd_sc_hd__dfrtp_1
X_9416_ clknet_leaf_10_csclk _0645_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][0]\ sky130_fd_sc_hd__dfstp_1
X_9417_ clknet_leaf_10_csclk _0646_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][1]\ sky130_fd_sc_hd__dfstp_1
X_9418_ clknet_leaf_9_csclk _0647_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][2]\ sky130_fd_sc_hd__dfrtp_1
X_9419_ clknet_leaf_10_csclk _0648_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][3]\ sky130_fd_sc_hd__dfrtp_2
X_9420_ clknet_leaf_10_csclk _0649_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][4]\ sky130_fd_sc_hd__dfrtp_1
X_9421_ clknet_leaf_10_csclk _0650_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][5]\ sky130_fd_sc_hd__dfrtp_2
X_9422_ clknet_leaf_10_csclk _0651_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][6]\ sky130_fd_sc_hd__dfrtp_1
X_9423_ clknet_leaf_10_csclk _0652_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][7]\ sky130_fd_sc_hd__dfrtp_1
X_9424_ clknet_leaf_12_csclk _0653_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][0]\ sky130_fd_sc_hd__dfstp_1
X_9425_ clknet_leaf_11_csclk _0654_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][1]\ sky130_fd_sc_hd__dfstp_1
X_9426_ clknet_leaf_11_csclk _0655_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][2]\ sky130_fd_sc_hd__dfrtp_1
X_9427_ clknet_leaf_11_csclk _0656_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][3]\ sky130_fd_sc_hd__dfrtp_1
X_9428_ clknet_leaf_17_csclk _0657_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][4]\ sky130_fd_sc_hd__dfrtp_1
X_9429_ clknet_leaf_17_csclk _0658_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][5]\ sky130_fd_sc_hd__dfrtp_1
X_9430_ clknet_leaf_17_csclk _0659_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][6]\ sky130_fd_sc_hd__dfrtp_1
X_9431_ clknet_leaf_17_csclk _0660_ net371 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[20][7]\ sky130_fd_sc_hd__dfrtp_1
X_9432_ clknet_leaf_6_csclk _0661_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][8]\ sky130_fd_sc_hd__dfrtp_1
X_9433_ clknet_leaf_6_csclk _0662_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][9]\ sky130_fd_sc_hd__dfrtp_1
X_9434_ clknet_leaf_6_csclk _0663_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][10]\ sky130_fd_sc_hd__dfstp_1
X_9435_ clknet_leaf_6_csclk _0664_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][11]\ sky130_fd_sc_hd__dfrtp_1
X_9436_ clknet_leaf_6_csclk _0665_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[32][12]\ sky130_fd_sc_hd__dfrtp_1
X_9437_ clknet_leaf_2_csclk _0666_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][8]\ sky130_fd_sc_hd__dfrtp_1
X_9438_ clknet_leaf_2_csclk _0667_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][9]\ sky130_fd_sc_hd__dfrtp_1
X_9439_ clknet_leaf_6_csclk _0668_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][10]\ sky130_fd_sc_hd__dfstp_1
X_9440_ clknet_leaf_6_csclk _0669_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][11]\ sky130_fd_sc_hd__dfrtp_1
X_9441_ clknet_leaf_2_csclk _0670_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][12]\ sky130_fd_sc_hd__dfrtp_1
X_9442_ clknet_leaf_36_csclk _0671_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][0]\ sky130_fd_sc_hd__dfstp_1
X_9443_ clknet_leaf_36_csclk _0672_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][1]\ sky130_fd_sc_hd__dfstp_1
X_9444_ clknet_leaf_40_csclk _0673_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][2]\ sky130_fd_sc_hd__dfrtp_1
X_9445_ clknet_leaf_36_csclk _0674_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][3]\ sky130_fd_sc_hd__dfrtp_4
X_9446_ clknet_leaf_36_csclk _0675_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][4]\ sky130_fd_sc_hd__dfrtp_1
X_9447_ clknet_leaf_36_csclk _0676_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][5]\ sky130_fd_sc_hd__dfrtp_1
X_9448_ clknet_leaf_40_csclk _0677_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][6]\ sky130_fd_sc_hd__dfrtp_1
X_9449_ clknet_leaf_40_csclk _0678_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][7]\ sky130_fd_sc_hd__dfrtp_1
X_9450_ clknet_leaf_18_csclk _0679_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][0]\ sky130_fd_sc_hd__dfstp_1
X_9451_ clknet_leaf_18_csclk _0680_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][1]\ sky130_fd_sc_hd__dfstp_1
X_9452_ clknet_leaf_18_csclk _0681_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][2]\ sky130_fd_sc_hd__dfrtp_1
X_9453_ clknet_leaf_18_csclk _0682_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][3]\ sky130_fd_sc_hd__dfrtp_1
X_9454_ clknet_leaf_18_csclk _0683_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][4]\ sky130_fd_sc_hd__dfrtp_1
X_9455_ clknet_leaf_18_csclk _0684_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][5]\ sky130_fd_sc_hd__dfrtp_1
X_9456_ clknet_leaf_19_csclk _0685_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][6]\ sky130_fd_sc_hd__dfrtp_1
X_9457_ clknet_leaf_18_csclk _0686_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[21][7]\ sky130_fd_sc_hd__dfrtp_1
X_9458_ clknet_leaf_5_csclk _0687_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][8]\ sky130_fd_sc_hd__dfrtp_1
X_9459_ clknet_leaf_13_csclk _0688_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][9]\ sky130_fd_sc_hd__dfrtp_1
X_9460_ clknet_leaf_13_csclk _0689_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][10]\ sky130_fd_sc_hd__dfstp_1
X_9461_ clknet_leaf_5_csclk _0690_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][11]\ sky130_fd_sc_hd__dfrtp_1
X_9462_ clknet_leaf_13_csclk _0691_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[31][12]\ sky130_fd_sc_hd__dfrtp_1
X_9463_ clknet_leaf_2_csclk _0692_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][8]\ sky130_fd_sc_hd__dfrtp_1
X_9464_ clknet_leaf_2_csclk _0693_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][9]\ sky130_fd_sc_hd__dfrtp_1
X_9465_ clknet_leaf_2_csclk _0694_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][10]\ sky130_fd_sc_hd__dfstp_1
X_9466_ clknet_leaf_2_csclk _0695_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][11]\ sky130_fd_sc_hd__dfrtp_1
X_9467_ clknet_leaf_2_csclk _0696_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][12]\ sky130_fd_sc_hd__dfrtp_1
X_9468_ clknet_leaf_12_csclk _0697_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][0]\ sky130_fd_sc_hd__dfstp_1
X_9469_ clknet_leaf_10_csclk _0698_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][1]\ sky130_fd_sc_hd__dfstp_1
X_9470_ clknet_leaf_9_csclk _0699_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][2]\ sky130_fd_sc_hd__dfrtp_1
X_9471_ clknet_leaf_9_csclk _0700_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][3]\ sky130_fd_sc_hd__dfrtp_4
X_9472_ clknet_leaf_10_csclk _0701_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][4]\ sky130_fd_sc_hd__dfrtp_1
X_9473_ clknet_leaf_9_csclk _0702_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][5]\ sky130_fd_sc_hd__dfrtp_2
X_9474_ clknet_leaf_9_csclk _0703_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][6]\ sky130_fd_sc_hd__dfrtp_1
X_9475_ clknet_leaf_9_csclk _0704_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][7]\ sky130_fd_sc_hd__dfrtp_1
X_9476_ clknet_leaf_11_csclk _0705_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][0]\ sky130_fd_sc_hd__dfstp_1
X_9477_ clknet_leaf_11_csclk _0706_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][1]\ sky130_fd_sc_hd__dfstp_1
X_9478_ clknet_leaf_18_csclk _0707_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][2]\ sky130_fd_sc_hd__dfrtp_1
X_9479_ clknet_leaf_10_csclk _0708_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][3]\ sky130_fd_sc_hd__dfrtp_4
X_9480_ clknet_leaf_11_csclk _0709_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][4]\ sky130_fd_sc_hd__dfrtp_1
X_9481_ clknet_leaf_11_csclk _0710_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][5]\ sky130_fd_sc_hd__dfrtp_1
X_9482_ clknet_leaf_18_csclk _0711_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][6]\ sky130_fd_sc_hd__dfrtp_1
X_9483_ clknet_leaf_18_csclk _0712_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[22][7]\ sky130_fd_sc_hd__dfrtp_1
X_9484_ clknet_leaf_45_csclk _0713_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][8]\ sky130_fd_sc_hd__dfrtp_1
X_9485_ clknet_leaf_48_csclk _0714_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][9]\ sky130_fd_sc_hd__dfrtp_1
X_9486_ clknet_leaf_45_csclk _0715_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][10]\ sky130_fd_sc_hd__dfstp_1
X_9487_ clknet_leaf_45_csclk _0716_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][11]\ sky130_fd_sc_hd__dfrtp_1
X_9488_ clknet_leaf_45_csclk _0717_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[30][12]\ sky130_fd_sc_hd__dfrtp_1
X_9489_ clknet_leaf_1_csclk _0718_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][8]\ sky130_fd_sc_hd__dfrtp_1
X_9490_ clknet_leaf_0_csclk _0719_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][9]\ sky130_fd_sc_hd__dfrtp_1
X_9491_ clknet_leaf_1_csclk _0720_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][10]\ sky130_fd_sc_hd__dfstp_1
X_9492_ clknet_leaf_0_csclk _0721_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][11]\ sky130_fd_sc_hd__dfrtp_1
X_9493_ clknet_leaf_1_csclk _0722_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][12]\ sky130_fd_sc_hd__dfrtp_1
X_9494_ clknet_leaf_14_csclk _0723_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][0]\ sky130_fd_sc_hd__dfstp_1
X_9495_ clknet_leaf_14_csclk _0724_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][1]\ sky130_fd_sc_hd__dfstp_1
X_9496_ clknet_leaf_13_csclk _0725_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][2]\ sky130_fd_sc_hd__dfrtp_1
X_9497_ clknet_leaf_15_csclk _0726_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][3]\ sky130_fd_sc_hd__dfrtp_4
X_9498_ clknet_leaf_14_csclk _0727_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][4]\ sky130_fd_sc_hd__dfrtp_1
X_9499_ clknet_leaf_15_csclk _0728_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][5]\ sky130_fd_sc_hd__dfrtp_1
X_9500_ clknet_leaf_15_csclk _0729_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][6]\ sky130_fd_sc_hd__dfrtp_1
X_9501_ clknet_leaf_15_csclk _0730_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][7]\ sky130_fd_sc_hd__dfrtp_1
X_9502_ clknet_leaf_11_csclk _0731_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][0]\ sky130_fd_sc_hd__dfstp_1
X_9503_ clknet_leaf_11_csclk _0732_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][1]\ sky130_fd_sc_hd__dfstp_1
X_9504_ clknet_leaf_17_csclk _0733_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][2]\ sky130_fd_sc_hd__dfrtp_1
X_9505_ clknet_leaf_11_csclk _0734_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][3]\ sky130_fd_sc_hd__dfrtp_1
X_9506_ clknet_leaf_11_csclk _0735_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][4]\ sky130_fd_sc_hd__dfrtp_1
X_9507_ clknet_leaf_19_csclk _0736_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][5]\ sky130_fd_sc_hd__dfrtp_1
X_9508_ clknet_leaf_17_csclk _0737_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][6]\ sky130_fd_sc_hd__dfrtp_1
X_9509_ clknet_leaf_19_csclk _0738_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[23][7]\ sky130_fd_sc_hd__dfrtp_1
X_9510_ clknet_leaf_2_csclk _0739_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][8]\ sky130_fd_sc_hd__dfrtp_1
X_9511_ clknet_leaf_2_csclk _0740_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][9]\ sky130_fd_sc_hd__dfrtp_1
X_9512_ clknet_leaf_2_csclk _0741_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][10]\ sky130_fd_sc_hd__dfstp_1
X_9513_ clknet_leaf_2_csclk _0742_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][11]\ sky130_fd_sc_hd__dfrtp_1
X_9514_ clknet_leaf_2_csclk _0743_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[29][12]\ sky130_fd_sc_hd__dfrtp_1
X_9515_ clknet_leaf_0_csclk _0744_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][8]\ sky130_fd_sc_hd__dfrtp_1
X_9516_ clknet_leaf_3_csclk _0745_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][9]\ sky130_fd_sc_hd__dfrtp_1
X_9517_ clknet_leaf_0_csclk _0746_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][10]\ sky130_fd_sc_hd__dfstp_1
X_9518_ clknet_leaf_0_csclk _0747_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][11]\ sky130_fd_sc_hd__dfrtp_1
X_9519_ clknet_leaf_3_csclk _0748_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][12]\ sky130_fd_sc_hd__dfrtp_1
X_9520_ clknet_leaf_11_csclk _0749_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][0]\ sky130_fd_sc_hd__dfstp_1
X_9521_ clknet_leaf_10_csclk _0750_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][1]\ sky130_fd_sc_hd__dfstp_1
X_9522_ clknet_leaf_11_csclk _0751_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][2]\ sky130_fd_sc_hd__dfrtp_1
X_9523_ clknet_leaf_10_csclk _0752_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][3]\ sky130_fd_sc_hd__dfrtp_2
X_9524_ clknet_leaf_11_csclk _0753_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][4]\ sky130_fd_sc_hd__dfrtp_1
X_9525_ clknet_leaf_10_csclk _0754_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][5]\ sky130_fd_sc_hd__dfrtp_1
X_9526_ clknet_leaf_11_csclk _0755_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][6]\ sky130_fd_sc_hd__dfrtp_1
X_9527_ clknet_leaf_11_csclk _0756_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][7]\ sky130_fd_sc_hd__dfrtp_1
X_9528_ clknet_leaf_12_csclk _0757_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][0]\ sky130_fd_sc_hd__dfstp_1
X_9529_ clknet_leaf_14_csclk _0758_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][1]\ sky130_fd_sc_hd__dfstp_1
X_9530_ clknet_leaf_13_csclk _0759_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][2]\ sky130_fd_sc_hd__dfrtp_1
X_9531_ clknet_leaf_12_csclk _0760_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][3]\ sky130_fd_sc_hd__dfrtp_4
X_9532_ clknet_leaf_13_csclk _0761_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][4]\ sky130_fd_sc_hd__dfrtp_1
X_9533_ clknet_leaf_12_csclk _0762_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][5]\ sky130_fd_sc_hd__dfrtp_1
X_9534_ clknet_leaf_14_csclk _0763_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][6]\ sky130_fd_sc_hd__dfrtp_1
X_9535_ clknet_leaf_12_csclk _0764_ net372 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[24][7]\ sky130_fd_sc_hd__dfrtp_1
X_9536_ clknet_leaf_51_csclk _0765_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][8]\ sky130_fd_sc_hd__dfrtp_1
X_9537_ clknet_leaf_51_csclk _0766_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][9]\ sky130_fd_sc_hd__dfrtp_1
X_9538_ clknet_leaf_51_csclk _0767_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][10]\ sky130_fd_sc_hd__dfstp_1
X_9539_ clknet_leaf_51_csclk _0768_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][11]\ sky130_fd_sc_hd__dfrtp_1
X_9540_ clknet_leaf_51_csclk _0769_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[28][12]\ sky130_fd_sc_hd__dfrtp_1
X_9541_ clknet_leaf_0_csclk _0770_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][8]\ sky130_fd_sc_hd__dfrtp_1
X_9542_ clknet_leaf_0_csclk _0771_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][9]\ sky130_fd_sc_hd__dfrtp_1
X_9543_ clknet_leaf_51_csclk _0772_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][10]\ sky130_fd_sc_hd__dfstp_1
X_9544_ clknet_leaf_51_csclk _0773_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][11]\ sky130_fd_sc_hd__dfrtp_1
X_9545_ clknet_leaf_0_csclk _0774_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][12]\ sky130_fd_sc_hd__dfrtp_1
X_9546_ clknet_leaf_38_csclk _0775_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][0]\ sky130_fd_sc_hd__dfstp_1
X_9547_ clknet_leaf_37_csclk _0776_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][1]\ sky130_fd_sc_hd__dfstp_1
X_9548_ clknet_leaf_37_csclk _0777_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][2]\ sky130_fd_sc_hd__dfrtp_1
X_9549_ clknet_leaf_37_csclk _0778_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][3]\ sky130_fd_sc_hd__dfrtp_2
X_9550_ clknet_leaf_39_csclk _0779_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][4]\ sky130_fd_sc_hd__dfrtp_1
X_9551_ clknet_leaf_37_csclk _0780_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][5]\ sky130_fd_sc_hd__dfrtp_1
X_9552_ clknet_leaf_37_csclk _0781_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][6]\ sky130_fd_sc_hd__dfrtp_1
X_9553_ clknet_leaf_37_csclk _0782_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][7]\ sky130_fd_sc_hd__dfrtp_1
X_9554_ clknet_leaf_44_csclk _0783_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][8]\ sky130_fd_sc_hd__dfrtp_1
X_9555_ clknet_leaf_43_csclk _0784_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][9]\ sky130_fd_sc_hd__dfrtp_1
X_9556_ clknet_leaf_45_csclk _0785_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][10]\ sky130_fd_sc_hd__dfstp_1
X_9557_ clknet_leaf_44_csclk _0786_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][11]\ sky130_fd_sc_hd__dfrtp_1
X_9558_ clknet_leaf_43_csclk _0787_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[27][12]\ sky130_fd_sc_hd__dfrtp_1
X_9559_ clknet_leaf_47_csclk _0788_ net375 VGND VGND VPWR 
+ VPWR
+ irq_1_inputsrc sky130_fd_sc_hd__dfrtp_1
X_9560_ clknet_leaf_47_csclk _0789_ net375 VGND VGND VPWR 
+ VPWR
+ irq_2_inputsrc sky130_fd_sc_hd__dfrtp_1
X_9561_ clknet_leaf_24_csclk _0790_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[16]\ sky130_fd_sc_hd__dfrtp_1
X_9562_ clknet_leaf_23_csclk _0791_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[17]\ sky130_fd_sc_hd__dfrtp_1
X_9563_ clknet_leaf_23_csclk _0792_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[18]\ sky130_fd_sc_hd__dfrtp_1
X_9564_ clknet_leaf_23_csclk _0793_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[19]\ sky130_fd_sc_hd__dfrtp_1
X_9565_ clknet_leaf_23_csclk _0794_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[20]\ sky130_fd_sc_hd__dfrtp_4
X_9566_ clknet_leaf_23_csclk _0795_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[21]\ sky130_fd_sc_hd__dfrtp_2
X_9567_ clknet_leaf_23_csclk _0796_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[22]\ sky130_fd_sc_hd__dfrtp_2
X_9568_ clknet_leaf_23_csclk _0797_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[23]\ sky130_fd_sc_hd__dfrtp_2
X_9569_ clknet_2_0_0_mgmt_gpio_in[4] _0798_ _0235_ VGND VGND VPWR 
+ VPWR
+ \hkspi.rdstb\ sky130_fd_sc_hd__dfrtp_2
X_9570_ clknet_leaf_26_csclk _0799_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[8]\ sky130_fd_sc_hd__dfrtp_2
X_9571_ clknet_leaf_26_csclk _0800_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[9]\ sky130_fd_sc_hd__dfrtp_1
X_9572_ clknet_leaf_24_csclk _0801_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[10]\ sky130_fd_sc_hd__dfrtp_2
X_9573_ clknet_leaf_26_csclk _0802_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[11]\ sky130_fd_sc_hd__dfrtp_1
X_9574_ clknet_leaf_24_csclk _0803_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[12]\ sky130_fd_sc_hd__dfrtp_1
X_9575_ clknet_leaf_26_csclk _0804_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[13]\ sky130_fd_sc_hd__dfrtp_1
X_9576_ clknet_leaf_24_csclk _0805_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[14]\ sky130_fd_sc_hd__dfrtp_1
X_9577_ clknet_leaf_24_csclk _0806_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[15]\ sky130_fd_sc_hd__dfrtp_1
X_9578_ clknet_leaf_33_csclk _0807_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[0]\ sky130_fd_sc_hd__dfrtp_1
X_9579_ clknet_leaf_33_csclk _0808_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[1]\ sky130_fd_sc_hd__dfrtp_4
X_9580_ clknet_leaf_34_csclk _0809_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[2]\ sky130_fd_sc_hd__dfrtp_1
X_9581_ clknet_leaf_34_csclk _0810_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[3]\ sky130_fd_sc_hd__dfrtp_1
X_9582_ clknet_leaf_33_csclk _0811_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[4]\ sky130_fd_sc_hd__dfrtp_1
X_9583_ clknet_leaf_33_csclk _0812_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[5]\ sky130_fd_sc_hd__dfrtp_1
X_9584_ clknet_leaf_33_csclk _0813_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[6]\ sky130_fd_sc_hd__dfrtp_1
X_9585_ clknet_leaf_33_csclk _0814_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[7]\ sky130_fd_sc_hd__dfrtp_2
X_9586_ clknet_2_0_0_mgmt_gpio_in[4] _0815_ _0236_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pass_thru_mgmt\ sky130_fd_sc_hd__dfrtp_4
X_9587_ clknet_3_6_0_wb_clk_i _0816_ net196 VGND VGND VPWR 
+ VPWR
+ wbbd_busy sky130_fd_sc_hd__dfrtp_4
X_9588_ clknet_leaf_22_csclk _0817_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[32]\ sky130_fd_sc_hd__dfrtp_1
X_9589_ clknet_leaf_23_csclk _0818_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[33]\ sky130_fd_sc_hd__dfrtp_1
X_9590_ clknet_leaf_22_csclk _0819_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[34]\ sky130_fd_sc_hd__dfrtp_1
X_9591_ clknet_leaf_22_csclk _0820_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[35]\ sky130_fd_sc_hd__dfrtp_1
X_9592_ clknet_leaf_23_csclk _0821_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[36]\ sky130_fd_sc_hd__dfrtp_1
X_9593_ clknet_leaf_22_csclk _0822_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[37]\ sky130_fd_sc_hd__dfrtp_1
X_9594_ clknet_leaf_20_csclk _0823_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[24]\ sky130_fd_sc_hd__dfrtp_1
X_9595_ clknet_leaf_20_csclk _0824_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[25]\ sky130_fd_sc_hd__dfrtp_1
X_9596_ clknet_leaf_20_csclk _0825_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[26]\ sky130_fd_sc_hd__dfrtp_1
X_9597_ clknet_leaf_22_csclk _0826_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[27]\ sky130_fd_sc_hd__dfrtp_1
X_9598_ clknet_leaf_22_csclk _0827_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[28]\ sky130_fd_sc_hd__dfrtp_1
X_9599_ clknet_leaf_22_csclk _0828_ net372 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[29]\ sky130_fd_sc_hd__dfrtp_1
X_9600_ clknet_leaf_22_csclk _0829_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[30]\ sky130_fd_sc_hd__dfrtp_1
X_9601_ clknet_leaf_22_csclk _0830_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data[31]\ sky130_fd_sc_hd__dfrtp_1
X_9602_ clknet_leaf_23_csclk _0831_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[16]\ sky130_fd_sc_hd__dfrtp_1
X_9603_ clknet_leaf_23_csclk _0832_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[17]\ sky130_fd_sc_hd__dfrtp_1
X_9604_ clknet_leaf_23_csclk _0833_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[18]\ sky130_fd_sc_hd__dfrtp_1
X_9605_ clknet_leaf_23_csclk _0834_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[19]\ sky130_fd_sc_hd__dfrtp_1
X_9606_ clknet_leaf_23_csclk _0835_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[20]\ sky130_fd_sc_hd__dfrtp_1
X_9607_ clknet_leaf_23_csclk _0836_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[21]\ sky130_fd_sc_hd__dfrtp_1
X_9608_ clknet_leaf_23_csclk _0837_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[22]\ sky130_fd_sc_hd__dfrtp_1
X_9609_ clknet_leaf_23_csclk _0838_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[23]\ sky130_fd_sc_hd__dfrtp_1
X_9610_ clknet_leaf_26_csclk _0839_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[8]\ sky130_fd_sc_hd__dfrtp_1
X_9611_ clknet_leaf_26_csclk _0840_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[9]\ sky130_fd_sc_hd__dfrtp_1
X_9612_ clknet_leaf_24_csclk _0841_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[10]\ sky130_fd_sc_hd__dfrtp_1
X_9613_ clknet_leaf_26_csclk _0842_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[11]\ sky130_fd_sc_hd__dfrtp_1
X_9614_ clknet_leaf_24_csclk _0843_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[12]\ sky130_fd_sc_hd__dfrtp_1
X_9615_ clknet_leaf_24_csclk _0844_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[13]\ sky130_fd_sc_hd__dfrtp_1
X_9616_ clknet_leaf_24_csclk _0845_ net369 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[14]\ sky130_fd_sc_hd__dfrtp_1
X_9617_ clknet_leaf_23_csclk _0846_ net371 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[15]\ sky130_fd_sc_hd__dfrtp_1
X_9618_ clknet_leaf_33_csclk _0847_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[0]\ sky130_fd_sc_hd__dfrtp_1
X_9619_ clknet_leaf_33_csclk _0848_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[1]\ sky130_fd_sc_hd__dfrtp_1
X_9620_ clknet_leaf_34_csclk _0849_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[2]\ sky130_fd_sc_hd__dfrtp_1
X_9621_ clknet_leaf_33_csclk _0850_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[3]\ sky130_fd_sc_hd__dfrtp_1
X_9622_ clknet_leaf_33_csclk _0851_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[4]\ sky130_fd_sc_hd__dfrtp_1
X_9623_ clknet_leaf_33_csclk _0852_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[5]\ sky130_fd_sc_hd__dfrtp_1
X_9624_ clknet_leaf_33_csclk _0853_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[6]\ sky130_fd_sc_hd__dfrtp_1
X_9625_ clknet_leaf_33_csclk _0854_ net376 VGND VGND VPWR 
+ VPWR
+ \mgmt_gpio_data_buf[7]\ sky130_fd_sc_hd__dfrtp_1
X_9626_ clknet_2_0_0_mgmt_gpio_in[4] _0855_ _0237_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pass_thru_mgmt_delay\ sky130_fd_sc_hd__dfrtp_4
X_9627_ clknet_leaf_38_csclk _0856_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][8]\ sky130_fd_sc_hd__dfrtp_1
X_9628_ clknet_leaf_37_csclk _0857_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][9]\ sky130_fd_sc_hd__dfrtp_1
X_9629_ clknet_leaf_38_csclk _0858_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][10]\ sky130_fd_sc_hd__dfrtp_2
X_9630_ clknet_leaf_37_csclk _0859_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][11]\ sky130_fd_sc_hd__dfstp_1
X_9631_ clknet_leaf_38_csclk _0860_ net377 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][12]\ sky130_fd_sc_hd__dfstp_1
X_9632_ clknet_leaf_37_csclk _0861_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][0]\ sky130_fd_sc_hd__dfstp_1
X_9633_ clknet_leaf_37_csclk _0862_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][1]\ sky130_fd_sc_hd__dfstp_1
X_9634_ clknet_leaf_39_csclk _0863_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][2]\ sky130_fd_sc_hd__dfrtp_1
X_9635_ clknet_leaf_36_csclk _0864_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][3]\ sky130_fd_sc_hd__dfrtp_1
X_9636_ clknet_leaf_37_csclk _0865_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][4]\ sky130_fd_sc_hd__dfrtp_1
X_9637_ clknet_leaf_36_csclk _0866_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][5]\ sky130_fd_sc_hd__dfrtp_1
X_9638_ clknet_leaf_37_csclk _0867_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][6]\ sky130_fd_sc_hd__dfrtp_1
X_9639_ clknet_leaf_37_csclk _0868_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[0][7]\ sky130_fd_sc_hd__dfrtp_1
X_9640_ clknet_3_6_0_wb_clk_i _0869_ net196 VGND VGND VPWR 
+ VPWR
+ wbbd_sck sky130_fd_sc_hd__dfrtp_2
X_9641_ clknet_leaf_48_csclk _0870_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][8]\ sky130_fd_sc_hd__dfrtp_1
X_9642_ clknet_leaf_47_csclk _0871_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][9]\ sky130_fd_sc_hd__dfrtp_1
X_9643_ clknet_leaf_47_csclk _0872_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][10]\ sky130_fd_sc_hd__dfrtp_1
X_9644_ clknet_leaf_47_csclk _0873_ net375 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][11]\ sky130_fd_sc_hd__dfstp_1
X_9645_ clknet_leaf_48_csclk _0874_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][12]\ sky130_fd_sc_hd__dfstp_1
X_9646_ clknet_leaf_25_csclk _0875_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][0]\ sky130_fd_sc_hd__dfstp_1
X_9647_ clknet_leaf_25_csclk _0876_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][1]\ sky130_fd_sc_hd__dfstp_1
X_9648_ clknet_leaf_25_csclk _0877_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][2]\ sky130_fd_sc_hd__dfrtp_1
X_9649_ clknet_leaf_25_csclk _0878_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][3]\ sky130_fd_sc_hd__dfrtp_1
X_9650_ clknet_leaf_29_csclk _0879_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][4]\ sky130_fd_sc_hd__dfrtp_1
X_9651_ clknet_leaf_29_csclk _0880_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][5]\ sky130_fd_sc_hd__dfrtp_1
X_9652_ clknet_leaf_25_csclk _0881_ net373 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][6]\ sky130_fd_sc_hd__dfrtp_1
X_9653_ clknet_leaf_29_csclk _0882_ net369 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[1][7]\ sky130_fd_sc_hd__dfrtp_1
X_9654_ clknet_leaf_41_csclk _0883_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][8]\ sky130_fd_sc_hd__dfrtp_1
X_9655_ clknet_leaf_39_csclk _0884_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][9]\ sky130_fd_sc_hd__dfrtp_1
X_9656_ clknet_leaf_41_csclk _0885_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][10]\ sky130_fd_sc_hd__dfstp_1
X_9657_ clknet_leaf_41_csclk _0886_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][11]\ sky130_fd_sc_hd__dfrtp_1
X_9658_ clknet_leaf_41_csclk _0887_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][12]\ sky130_fd_sc_hd__dfrtp_1
X_9659_ clknet_3_6_0_wb_clk_i _0888_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[0]\ sky130_fd_sc_hd__dfrtp_1
X_9660_ clknet_3_7_0_wb_clk_i _0889_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[1]\ sky130_fd_sc_hd__dfrtp_1
X_9661_ clknet_3_7_0_wb_clk_i _0890_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[2]\ sky130_fd_sc_hd__dfrtp_1
X_9662_ clknet_3_7_0_wb_clk_i _0891_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[3]\ sky130_fd_sc_hd__dfrtp_1
X_9663_ clknet_3_7_0_wb_clk_i _0892_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[4]\ sky130_fd_sc_hd__dfrtp_1
X_9664_ clknet_3_7_0_wb_clk_i _0893_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[5]\ sky130_fd_sc_hd__dfrtp_1
X_9665_ clknet_3_6_0_wb_clk_i _0894_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[6]\ sky130_fd_sc_hd__dfrtp_1
X_9666_ clknet_3_6_0_wb_clk_i _0895_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_data[7]\ sky130_fd_sc_hd__dfrtp_1
X_9667_ clknet_leaf_33_csclk _0896_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][0]\ sky130_fd_sc_hd__dfstp_1
X_9668_ clknet_leaf_33_csclk _0897_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][1]\ sky130_fd_sc_hd__dfstp_1
X_9669_ clknet_leaf_33_csclk _0898_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][2]\ sky130_fd_sc_hd__dfrtp_1
X_9670_ clknet_leaf_33_csclk _0899_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][3]\ sky130_fd_sc_hd__dfrtp_1
X_9671_ clknet_leaf_33_csclk _0900_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][4]\ sky130_fd_sc_hd__dfrtp_1
X_9672_ clknet_leaf_32_csclk _0901_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][5]\ sky130_fd_sc_hd__dfrtp_1
X_9673_ clknet_leaf_33_csclk _0902_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][6]\ sky130_fd_sc_hd__dfrtp_1
X_9674_ clknet_leaf_33_csclk _0903_ net376 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[2][7]\ sky130_fd_sc_hd__dfrtp_1
X_9675_ clknet_3_1_0_wb_clk_i _0904_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[0]\ sky130_fd_sc_hd__dfrtp_1
X_9676_ clknet_3_1_0_wb_clk_i _0905_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[1]\ sky130_fd_sc_hd__dfrtp_1
X_9677_ clknet_3_1_0_wb_clk_i _0906_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[2]\ sky130_fd_sc_hd__dfrtp_1
X_9678_ clknet_3_1_0_wb_clk_i _0907_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[3]\ sky130_fd_sc_hd__dfrtp_1
X_9679_ clknet_3_1_0_wb_clk_i _0908_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[4]\ sky130_fd_sc_hd__dfrtp_1
X_9680_ clknet_3_1_0_wb_clk_i _0909_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[5]\ sky130_fd_sc_hd__dfrtp_1
X_9681_ clknet_3_1_0_wb_clk_i _0910_ net196 VGND VGND VPWR 
+ VPWR
+ \wbbd_addr[6]\ sky130_fd_sc_hd__dfrtp_1
X_9682_ clknet_2_1_0_mgmt_gpio_in[4] _0911_ _0238_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pass_thru_user\ sky130_fd_sc_hd__dfrtp_4
X_9683_ clknet_leaf_10_csclk _0912_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][8]\ sky130_fd_sc_hd__dfrtp_1
X_9684_ clknet_leaf_10_csclk _0913_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][9]\ sky130_fd_sc_hd__dfrtp_1
X_9685_ clknet_leaf_9_csclk _0914_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][10]\ sky130_fd_sc_hd__dfstp_1
X_9686_ clknet_leaf_9_csclk _0915_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][11]\ sky130_fd_sc_hd__dfrtp_1
X_9687_ clknet_leaf_9_csclk _0916_ net374 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[3][12]\ sky130_fd_sc_hd__dfrtp_1
X_9688_ clknet_leaf_32_csclk _0917_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][0]\ sky130_fd_sc_hd__dfstp_1
X_9689_ clknet_leaf_32_csclk _0918_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][1]\ sky130_fd_sc_hd__dfstp_1
X_9690_ clknet_leaf_32_csclk _0919_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][2]\ sky130_fd_sc_hd__dfrtp_1
X_9691_ clknet_leaf_32_csclk _0920_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][3]\ sky130_fd_sc_hd__dfrtp_1
X_9692_ clknet_leaf_32_csclk _0921_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][4]\ sky130_fd_sc_hd__dfrtp_1
X_9693_ clknet_leaf_32_csclk _0922_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][5]\ sky130_fd_sc_hd__dfrtp_1
X_9694_ clknet_leaf_32_csclk _0923_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][6]\ sky130_fd_sc_hd__dfrtp_1
X_9695_ clknet_leaf_32_csclk _0924_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[5][7]\ sky130_fd_sc_hd__dfrtp_1
X_9696_ clknet_2_0_0_mgmt_gpio_in[4] _0925_ _0239_ VGND VGND VPWR 
+ VPWR
+ \hkspi.writemode\ sky130_fd_sc_hd__dfrtp_1
X_9697_ clknet_2_1_0_mgmt_gpio_in[4] _0926_ _0240_ VGND VGND VPWR 
+ VPWR
+ \hkspi.readmode\ sky130_fd_sc_hd__dfrtp_1
X_9698_ clknet_2_1_0_mgmt_gpio_in[4] _0927_ _0241_ VGND VGND VPWR 
+ VPWR
+ \hkspi.fixed[0]\ sky130_fd_sc_hd__dfrtp_4
X_9699_ clknet_2_1_0_mgmt_gpio_in[4] _0928_ _0242_ VGND VGND VPWR 
+ VPWR
+ \hkspi.fixed[1]\ sky130_fd_sc_hd__dfrtp_1
X_9700_ clknet_2_1_0_mgmt_gpio_in[4] _0929_ _0243_ VGND VGND VPWR 
+ VPWR
+ \hkspi.fixed[2]\ sky130_fd_sc_hd__dfrtp_1
X_9701_ clknet_2_3_0_mgmt_gpio_in[4] _0930_ _0244_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[1]\ sky130_fd_sc_hd__dfrtp_1
X_9702_ clknet_2_3_0_mgmt_gpio_in[4] _0931_ _0245_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[2]\ sky130_fd_sc_hd__dfrtp_1
X_9703_ clknet_2_3_0_mgmt_gpio_in[4] _0932_ _0246_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[3]\ sky130_fd_sc_hd__dfrtp_1
X_9704_ clknet_2_3_0_mgmt_gpio_in[4] _0933_ _0247_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[4]\ sky130_fd_sc_hd__dfrtp_1
X_9705_ clknet_2_3_0_mgmt_gpio_in[4] _0934_ _0248_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[5]\ sky130_fd_sc_hd__dfrtp_1
X_9706_ clknet_2_3_0_mgmt_gpio_in[4] _0935_ _0249_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[6]\ sky130_fd_sc_hd__dfrtp_1
X_9707_ clknet_2_3_0_mgmt_gpio_in[4] _0936_ _0250_ VGND VGND VPWR 
+ VPWR
+ \hkspi.odata[7]\ sky130_fd_sc_hd__dfrtp_1
X_9708_ clknet_2_1_0_mgmt_gpio_in[4] _0937_ _0251_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pre_pass_thru_mgmt\ sky130_fd_sc_hd__dfrtp_2
X_9709_ clknet_2_1_0_mgmt_gpio_in[4] _0938_ _0252_ VGND VGND VPWR 
+ VPWR
+ \hkspi.pre_pass_thru_user\ sky130_fd_sc_hd__dfrtp_1
X_9710_ clknet_2_1_0_mgmt_gpio_in[4] _0939_ _0253_ VGND VGND VPWR 
+ VPWR
+ \hkspi.wrstb\ sky130_fd_sc_hd__dfrtn_1
X_9711_ clknet_2_1_0_mgmt_gpio_in[4] _0940_ _0254_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[0]\ sky130_fd_sc_hd__dfrtn_1
X_9712_ clknet_2_2_0_mgmt_gpio_in[4] _0941_ _0255_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[1]\ sky130_fd_sc_hd__dfrtn_1
X_9713_ clknet_2_2_0_mgmt_gpio_in[4] _0942_ _0256_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[2]\ sky130_fd_sc_hd__dfrtn_1
X_9714_ clknet_2_2_0_mgmt_gpio_in[4] _0943_ _0257_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[3]\ sky130_fd_sc_hd__dfrtn_1
X_9715_ clknet_2_2_0_mgmt_gpio_in[4] _0944_ _0258_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[4]\ sky130_fd_sc_hd__dfrtn_1
X_9716_ clknet_2_2_0_mgmt_gpio_in[4] _0945_ _0259_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[5]\ sky130_fd_sc_hd__dfrtn_1
X_9717_ clknet_2_1_0_mgmt_gpio_in[4] net394 _0260_ VGND VGND VPWR 
+ VPWR
+ \hkspi.ldata[6]\ sky130_fd_sc_hd__dfrtn_1
X_9718_ clknet_2_0_0_mgmt_gpio_in[4] _0947_ _0261_ VGND VGND VPWR 
+ VPWR
+ \hkspi.SDO\ sky130_fd_sc_hd__dfrtn_1
X_9719_ clknet_leaf_50_csclk _0948_ net75 VGND VGND VPWR 
+ VPWR
+ net270 sky130_fd_sc_hd__dfrtp_1
X_9720_ clknet_leaf_50_csclk _0949_ net75 VGND VGND VPWR 
+ VPWR
+ net264 sky130_fd_sc_hd__dfstp_1
X_9721_ clknet_leaf_49_csclk _0950_ net377 VGND VGND VPWR 
+ VPWR
+ net265 sky130_fd_sc_hd__dfrtp_1
X_9722_ clknet_leaf_49_csclk _0951_ net75 VGND VGND VPWR 
+ VPWR
+ net266 sky130_fd_sc_hd__dfrtp_2
X_9723_ clknet_leaf_49_csclk _0952_ net377 VGND VGND VPWR 
+ VPWR
+ net267 sky130_fd_sc_hd__dfstp_1
X_9724_ clknet_leaf_49_csclk _0953_ net377 VGND VGND VPWR 
+ VPWR
+ net268 sky130_fd_sc_hd__dfrtp_1
X_9725_ clknet_leaf_49_csclk _0954_ net377 VGND VGND VPWR 
+ VPWR
+ net269 sky130_fd_sc_hd__dfrtp_1
X_9726_ clknet_leaf_49_csclk _0955_ net75 VGND VGND VPWR 
+ VPWR
+ net271 sky130_fd_sc_hd__dfrtp_2
X_9727_ clknet_leaf_49_csclk _0956_ net75 VGND VGND VPWR 
+ VPWR
+ net272 sky130_fd_sc_hd__dfstp_1
X_9728_ clknet_leaf_49_csclk _0957_ net75 VGND VGND VPWR 
+ VPWR
+ net273 sky130_fd_sc_hd__dfrtp_2
X_9729_ clknet_leaf_48_csclk _0958_ net377 VGND VGND VPWR 
+ VPWR
+ net260 sky130_fd_sc_hd__dfrtp_1
X_9730_ clknet_leaf_48_csclk _0959_ net75 VGND VGND VPWR 
+ VPWR
+ net261 sky130_fd_sc_hd__dfstp_2
X_9731_ clknet_leaf_48_csclk _0960_ net75 VGND VGND VPWR 
+ VPWR
+ net262 sky130_fd_sc_hd__dfrtp_1
X_9732_ clknet_leaf_48_csclk _0961_ net377 VGND VGND VPWR 
+ VPWR
+ net274 sky130_fd_sc_hd__dfstp_1
X_9733_ clknet_leaf_48_csclk _0962_ net377 VGND VGND VPWR 
+ VPWR
+ net285 sky130_fd_sc_hd__dfstp_1
X_9734_ clknet_leaf_48_csclk _0963_ net377 VGND VGND VPWR 
+ VPWR
+ net292 sky130_fd_sc_hd__dfstp_1
X_9735_ clknet_leaf_48_csclk _0964_ net377 VGND VGND VPWR 
+ VPWR
+ net293 sky130_fd_sc_hd__dfstp_1
X_9736_ clknet_leaf_48_csclk _0965_ net377 VGND VGND VPWR 
+ VPWR
+ net294 sky130_fd_sc_hd__dfstp_1
X_9737_ clknet_leaf_48_csclk _0966_ net377 VGND VGND VPWR 
+ VPWR
+ net295 sky130_fd_sc_hd__dfstp_1
X_9738_ clknet_leaf_48_csclk _0967_ net377 VGND VGND VPWR 
+ VPWR
+ net296 sky130_fd_sc_hd__dfstp_1
X_9739_ clknet_leaf_48_csclk _0968_ net377 VGND VGND VPWR 
+ VPWR
+ net297 sky130_fd_sc_hd__dfstp_1
X_9740_ clknet_leaf_45_csclk _0969_ net377 VGND VGND VPWR 
+ VPWR
+ net298 sky130_fd_sc_hd__dfstp_1
X_9741_ clknet_leaf_45_csclk _0970_ net377 VGND VGND VPWR 
+ VPWR
+ net299 sky130_fd_sc_hd__dfstp_1
X_9742_ clknet_leaf_45_csclk _0971_ net377 VGND VGND VPWR 
+ VPWR
+ net275 sky130_fd_sc_hd__dfstp_1
X_9743_ clknet_leaf_45_csclk _0972_ net377 VGND VGND VPWR 
+ VPWR
+ net276 sky130_fd_sc_hd__dfstp_1
X_9744_ clknet_leaf_45_csclk _0973_ net377 VGND VGND VPWR 
+ VPWR
+ net277 sky130_fd_sc_hd__dfrtp_1
X_9745_ clknet_leaf_45_csclk _0974_ net377 VGND VGND VPWR 
+ VPWR
+ net278 sky130_fd_sc_hd__dfstp_1
X_9746_ clknet_leaf_45_csclk _0975_ net377 VGND VGND VPWR 
+ VPWR
+ net279 sky130_fd_sc_hd__dfstp_1
X_9747_ clknet_leaf_45_csclk _0976_ net377 VGND VGND VPWR 
+ VPWR
+ net280 sky130_fd_sc_hd__dfstp_1
X_9748_ clknet_leaf_44_csclk _0977_ net377 VGND VGND VPWR 
+ VPWR
+ net281 sky130_fd_sc_hd__dfstp_1
X_9749_ clknet_leaf_45_csclk _0978_ net377 VGND VGND VPWR 
+ VPWR
+ net282 sky130_fd_sc_hd__dfstp_1
X_9750_ clknet_leaf_44_csclk _0979_ net377 VGND VGND VPWR 
+ VPWR
+ net283 sky130_fd_sc_hd__dfstp_1
X_9751_ clknet_leaf_44_csclk _0980_ net377 VGND VGND VPWR 
+ VPWR
+ net284 sky130_fd_sc_hd__dfstp_1
X_9752_ clknet_leaf_44_csclk _0981_ net377 VGND VGND VPWR 
+ VPWR
+ net286 sky130_fd_sc_hd__dfstp_1
X_9753_ clknet_leaf_44_csclk _0982_ net377 VGND VGND VPWR 
+ VPWR
+ net287 sky130_fd_sc_hd__dfstp_1
X_9754_ clknet_leaf_44_csclk _0983_ net377 VGND VGND VPWR 
+ VPWR
+ net288 sky130_fd_sc_hd__dfstp_1
X_9755_ clknet_leaf_44_csclk _0984_ net377 VGND VGND VPWR 
+ VPWR
+ net289 sky130_fd_sc_hd__dfstp_1
X_9756_ clknet_leaf_38_csclk _0985_ net377 VGND VGND VPWR 
+ VPWR
+ net290 sky130_fd_sc_hd__dfstp_1
X_9757_ clknet_leaf_38_csclk _0986_ net377 VGND VGND VPWR 
+ VPWR
+ net291 sky130_fd_sc_hd__dfstp_1
X_9758_ clknet_leaf_43_csclk _0987_ net75 VGND VGND VPWR 
+ VPWR
+ net263 sky130_fd_sc_hd__dfstp_1
X_9759_ clknet_3_6_0_wb_clk_i _0988_ net196 VGND VGND VPWR 
+ VPWR
+ wbbd_write sky130_fd_sc_hd__dfrtp_4
X_9760_ clknet_leaf_50_csclk _0989_ net75 VGND VGND VPWR 
+ VPWR
+ net324 sky130_fd_sc_hd__dfrtp_1
X_9761_ clknet_leaf_50_csclk _0990_ net75 VGND VGND VPWR 
+ VPWR
+ net325 sky130_fd_sc_hd__dfstp_2
X_9762_ clknet_leaf_50_csclk _0991_ net75 VGND VGND VPWR 
+ VPWR
+ net316 sky130_fd_sc_hd__dfrtp_4
X_9763_ clknet_leaf_50_csclk _0992_ net75 VGND VGND VPWR 
+ VPWR
+ net317 sky130_fd_sc_hd__dfrtp_2
X_9764_ clknet_leaf_50_csclk _0993_ net75 VGND VGND VPWR 
+ VPWR
+ net318 sky130_fd_sc_hd__dfrtp_4
X_9765_ clknet_leaf_51_csclk _0994_ net375 VGND VGND VPWR 
+ VPWR
+ net319 sky130_fd_sc_hd__dfrtp_4
X_9766_ clknet_leaf_49_csclk _0995_ net377 VGND VGND VPWR 
+ VPWR
+ net320 sky130_fd_sc_hd__dfrtp_2
X_9767_ clknet_leaf_49_csclk _0996_ net377 VGND VGND VPWR 
+ VPWR
+ net321 sky130_fd_sc_hd__dfrtp_2
X_9768_ clknet_leaf_51_csclk _0997_ net375 VGND VGND VPWR 
+ VPWR
+ net322 sky130_fd_sc_hd__dfrtp_4
X_9769_ clknet_leaf_49_csclk _0998_ net375 VGND VGND VPWR 
+ VPWR
+ net323 sky130_fd_sc_hd__dfrtp_4
X_9770_ clknet_leaf_50_csclk _0999_ net75 VGND VGND VPWR 
+ VPWR
+ reset_reg sky130_fd_sc_hd__dfrtp_1
X_9771_ clknet_leaf_3_csclk _1000_ net375 VGND VGND VPWR 
+ VPWR
+ net204 sky130_fd_sc_hd__dfrtp_2
X_9772_ clknet_leaf_35_csclk _1001_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_clock sky130_fd_sc_hd__dfrtp_2
X_9773_ clknet_leaf_46_csclk _1002_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][8]\ sky130_fd_sc_hd__dfrtp_1
X_9774_ clknet_leaf_48_csclk _1003_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][9]\ sky130_fd_sc_hd__dfrtp_1
X_9775_ clknet_leaf_46_csclk _1004_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][10]\ sky130_fd_sc_hd__dfstp_1
X_9776_ clknet_leaf_47_csclk _1005_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][11]\ sky130_fd_sc_hd__dfrtp_1
X_9777_ clknet_leaf_45_csclk _1006_ net75 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[26][12]\ sky130_fd_sc_hd__dfrtp_1
X_9778_ clknet_leaf_40_csclk _1007_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][0]\ sky130_fd_sc_hd__dfstp_1
X_9779_ clknet_leaf_41_csclk _1008_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][1]\ sky130_fd_sc_hd__dfstp_1
X_9780_ clknet_leaf_40_csclk _1009_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][2]\ sky130_fd_sc_hd__dfrtp_1
X_9781_ clknet_leaf_40_csclk _1010_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][3]\ sky130_fd_sc_hd__dfrtp_1
X_9782_ clknet_leaf_40_csclk _1011_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][4]\ sky130_fd_sc_hd__dfrtp_1
X_9783_ clknet_leaf_40_csclk _1012_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][5]\ sky130_fd_sc_hd__dfrtp_1
X_9784_ clknet_leaf_40_csclk _1013_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][6]\ sky130_fd_sc_hd__dfrtp_1
X_9785_ clknet_leaf_40_csclk _1014_ net370 VGND VGND VPWR 
+ VPWR
+ \gpio_configure[25][7]\ sky130_fd_sc_hd__dfrtp_1
X_9786_ clknet_leaf_24_csclk _1015_ net371 VGND VGND VPWR 
+ VPWR
+ clk2_output_dest sky130_fd_sc_hd__dfrtp_1
X_9787_ clknet_leaf_35_csclk _1016_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_enable sky130_fd_sc_hd__dfrtp_4
X_9788_ clknet_leaf_24_csclk _1017_ net369 VGND VGND VPWR 
+ VPWR
+ clk1_output_dest sky130_fd_sc_hd__dfrtp_2
X_9789_ clknet_leaf_5_csclk _1018_ net374 VGND VGND VPWR 
+ VPWR
+ hkspi_disable sky130_fd_sc_hd__dfrtp_1
X_9790_ clknet_leaf_35_csclk _1019_ net377 VGND VGND VPWR 
+ VPWR
+ serial_bb_data_2 sky130_fd_sc_hd__dfrtp_1
X_9791_ clknet_leaf_36_csclk _1020_ net376 VGND VGND VPWR 
+ VPWR
+ serial_xfer sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_csclk csclk VGND VGND VPWR VPWR clknet_0_csclk sky130_fd_sc_hd__clkbuf_16
X\clkbuf_0_mgmt_gpio_in[4]  mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0_wb_clk_i wb_clk_i VGND VGND VPWR VPWR clknet_0_wb_clk_i sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0_csclk clknet_0_csclk VGND VGND VPWR VPWR clknet_1_0_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_1_0_0_mgmt_gpio_in[4]  clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_1_0_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_0_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_1_csclk clknet_1_0_0_csclk VGND VGND VPWR VPWR clknet_1_0_1_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_1_0_1_mgmt_gpio_in[4]  clknet_1_0_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_1_0_1_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_1_wb_clk_i clknet_1_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_0_1_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_csclk clknet_0_csclk VGND VGND VPWR VPWR clknet_1_1_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_1_1_0_mgmt_gpio_in[4]  clknet_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_1_1_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_wb_clk_i clknet_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_1_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_1_csclk clknet_1_1_0_csclk VGND VGND VPWR VPWR clknet_1_1_1_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_1_1_1_mgmt_gpio_in[4]  clknet_1_1_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_1_1_1_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_1_wb_clk_i clknet_1_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_1_1_1_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_0_0_csclk clknet_1_0_1_csclk VGND VGND VPWR VPWR clknet_2_0_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_2_0_0_mgmt_gpio_in[4]  clknet_1_0_1_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_0_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_0_0_wb_clk_i clknet_1_0_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_0_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_csclk clknet_1_0_1_csclk VGND VGND VPWR VPWR clknet_2_1_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_2_1_0_mgmt_gpio_in[4]  clknet_1_0_1_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_1_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_1_0_wb_clk_i clknet_1_0_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_1_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_2_0_csclk clknet_1_1_1_csclk VGND VGND VPWR VPWR clknet_2_2_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_2_2_0_mgmt_gpio_in[4]  clknet_1_1_1_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_2_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_2_0_wb_clk_i clknet_1_1_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_2_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_3_0_csclk clknet_1_1_1_csclk VGND VGND VPWR VPWR clknet_2_3_0_csclk sky130_fd_sc_hd__clkbuf_2
X\clkbuf_2_3_0_mgmt_gpio_in[4]  clknet_1_1_1_mgmt_gpio_in[4] VGND VGND VPWR VPWR clknet_2_3_0_mgmt_gpio_in[4] sky130_fd_sc_hd__clkbuf_2
Xclkbuf_2_3_0_wb_clk_i clknet_1_1_1_wb_clk_i VGND VGND VPWR VPWR clknet_2_3_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_0_0_wb_clk_i clknet_2_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_0_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_1_0_wb_clk_i clknet_2_0_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_1_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_2_0_wb_clk_i clknet_2_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_2_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_3_0_wb_clk_i clknet_2_1_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_3_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_4_0_wb_clk_i clknet_2_2_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_4_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_5_0_wb_clk_i clknet_2_2_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_5_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_6_0_wb_clk_i clknet_2_3_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_6_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_3_7_0_wb_clk_i clknet_2_3_0_wb_clk_i VGND VGND VPWR VPWR clknet_3_7_0_wb_clk_i sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_0_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_10_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_10_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_11_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_11_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_12_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_12_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_13_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_13_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_14_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_14_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_15_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_15_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_16_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_16_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_17_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_17_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_18_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_18_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_19_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_19_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_1_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_1_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_20_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_20_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_21_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_21_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_22_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_22_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_23_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_23_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_24_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_24_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_25_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_25_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_26_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_26_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_27_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_27_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_28_csclk clknet_opt_6_0_csclk VGND VGND VPWR VPWR clknet_leaf_28_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_29_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_29_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_2_csclk clknet_opt_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_2_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_30_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_30_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_31_csclk clknet_opt_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_31_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_32_csclk clknet_opt_3_0_csclk VGND VGND VPWR VPWR clknet_leaf_32_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_33_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_33_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_34_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_34_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_35_csclk clknet_opt_4_0_csclk VGND VGND VPWR VPWR clknet_leaf_35_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_36_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_36_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_37_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_37_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_38_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_38_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_39_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_39_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_3_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_3_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_40_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_40_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_41_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_leaf_41_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_43_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_43_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_44_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_44_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_45_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_45_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_46_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_46_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_47_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_47_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_48_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_48_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_49_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_49_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_4_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_4_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_50_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_50_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_51_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_leaf_51_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_5_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_5_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_6_csclk clknet_opt_5_0_csclk VGND VGND VPWR VPWR clknet_leaf_6_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_7_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_7_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_8_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_8_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_leaf_9_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_leaf_9_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_1_0_csclk clknet_2_0_0_csclk VGND VGND VPWR VPWR clknet_opt_1_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_2_0_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_opt_2_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_3_0_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_opt_3_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_4_0_csclk clknet_2_1_0_csclk VGND VGND VPWR VPWR clknet_opt_4_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_5_0_csclk clknet_2_2_0_csclk VGND VGND VPWR VPWR clknet_opt_5_0_csclk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_opt_6_0_csclk clknet_2_3_0_csclk VGND VGND VPWR VPWR clknet_opt_6_0_csclk sky130_fd_sc_hd__clkbuf_16
Xhold1 \hkspi.ldata[5]\ VGND VGND VPWR VPWR net393 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2 _0946_ VGND VGND VPWR VPWR net394 sky130_fd_sc_hd__clkdlybuf4s25_1
Xinput1 debug_mode VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_4
Xinput10 mask_rev_in[15] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
Xinput100 sram_ro_data[16] VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
Xinput101 sram_ro_data[17] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xinput102 sram_ro_data[18] VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
Xinput103 sram_ro_data[19] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
Xinput104 sram_ro_data[1] VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
Xinput105 sram_ro_data[20] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput106 sram_ro_data[21] VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__clkbuf_1
Xinput107 sram_ro_data[22] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
Xinput108 sram_ro_data[23] VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__clkbuf_1
Xinput109 sram_ro_data[24] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__clkbuf_1
Xinput11 mask_rev_in[16] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
Xinput110 sram_ro_data[25] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__clkbuf_1
Xinput111 sram_ro_data[26] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
Xinput112 sram_ro_data[27] VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__clkbuf_1
Xinput113 sram_ro_data[28] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
Xinput114 sram_ro_data[29] VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__clkbuf_1
Xinput115 sram_ro_data[2] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__clkbuf_1
Xinput116 sram_ro_data[30] VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__clkbuf_1
Xinput117 sram_ro_data[31] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__clkbuf_1
Xinput118 sram_ro_data[3] VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__clkbuf_1
Xinput119 sram_ro_data[4] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__clkbuf_1
Xinput12 mask_rev_in[17] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
Xinput120 sram_ro_data[5] VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__clkbuf_1
Xinput121 sram_ro_data[6] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__clkbuf_1
Xinput122 sram_ro_data[7] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__clkbuf_1
Xinput123 sram_ro_data[8] VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__clkbuf_1
Xinput124 sram_ro_data[9] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__clkbuf_1
Xinput125 trap VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__buf_6
Xinput126 uart_enabled VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__buf_4
Xinput127 usr1_vcc_pwrgood VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__clkbuf_1
Xinput128 usr1_vdd_pwrgood VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__clkbuf_1
Xinput129 usr2_vcc_pwrgood VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__clkbuf_1
Xinput13 mask_rev_in[18] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput130 usr2_vdd_pwrgood VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__clkbuf_1
Xinput131 wb_adr_i[0] VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__clkbuf_4
Xinput132 wb_adr_i[10] VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__clkbuf_1
Xinput133 wb_adr_i[11] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__clkbuf_1
Xinput134 wb_adr_i[12] VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__clkbuf_1
Xinput135 wb_adr_i[13] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__clkbuf_1
Xinput136 wb_adr_i[14] VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__clkbuf_1
Xinput137 wb_adr_i[15] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__clkbuf_1
Xinput138 wb_adr_i[16] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__clkbuf_1
Xinput139 wb_adr_i[17] VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__clkbuf_1
Xinput14 mask_rev_in[19] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput140 wb_adr_i[18] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__clkbuf_1
Xinput141 wb_adr_i[19] VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_1
Xinput142 wb_adr_i[1] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_4
Xinput143 wb_adr_i[20] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__buf_2
Xinput144 wb_adr_i[21] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_2
Xinput145 wb_adr_i[22] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_1
Xinput146 wb_adr_i[23] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_1
Xinput147 wb_adr_i[24] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__clkbuf_1
Xinput148 wb_adr_i[25] VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_1
Xinput149 wb_adr_i[26] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__clkbuf_1
Xinput15 mask_rev_in[1] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xinput150 wb_adr_i[27] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_1
Xinput151 wb_adr_i[28] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_1
Xinput152 wb_adr_i[29] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_1
Xinput153 wb_adr_i[2] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__buf_4
Xinput154 wb_adr_i[30] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_1
Xinput155 wb_adr_i[31] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_1
Xinput156 wb_adr_i[3] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__buf_4
Xinput157 wb_adr_i[4] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__buf_4
Xinput158 wb_adr_i[5] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__buf_6
Xinput159 wb_adr_i[6] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__buf_4
Xinput16 mask_rev_in[20] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xinput160 wb_adr_i[7] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_6
Xinput161 wb_adr_i[8] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__clkbuf_1
Xinput162 wb_adr_i[9] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__clkbuf_1
Xinput163 wb_cyc_i VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput164 wb_dat_i[0] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_1
Xinput165 wb_dat_i[10] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_1
Xinput166 wb_dat_i[11] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_1
Xinput167 wb_dat_i[12] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_1
Xinput168 wb_dat_i[13] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_1
Xinput169 wb_dat_i[14] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_1
Xinput17 mask_rev_in[21] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
Xinput170 wb_dat_i[15] VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_1
Xinput171 wb_dat_i[16] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__clkbuf_1
Xinput172 wb_dat_i[17] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__clkbuf_1
Xinput173 wb_dat_i[18] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_1
Xinput174 wb_dat_i[19] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_1
Xinput175 wb_dat_i[1] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_1
Xinput176 wb_dat_i[20] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_1
Xinput177 wb_dat_i[21] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__clkbuf_1
Xinput178 wb_dat_i[22] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_1
Xinput179 wb_dat_i[23] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_1
Xinput18 mask_rev_in[22] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
Xinput180 wb_dat_i[24] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_1
Xinput181 wb_dat_i[25] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_1
Xinput182 wb_dat_i[26] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__clkbuf_1
Xinput183 wb_dat_i[27] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_1
Xinput184 wb_dat_i[28] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_1
Xinput185 wb_dat_i[29] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_1
Xinput186 wb_dat_i[2] VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_1
Xinput187 wb_dat_i[30] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_1
Xinput188 wb_dat_i[31] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_1
Xinput189 wb_dat_i[3] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_1
Xinput19 mask_rev_in[23] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
Xinput190 wb_dat_i[4] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_1
Xinput191 wb_dat_i[5] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_1
Xinput192 wb_dat_i[6] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_1
Xinput193 wb_dat_i[7] VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__clkbuf_1
Xinput194 wb_dat_i[8] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_1
Xinput195 wb_dat_i[9] VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__clkbuf_1
Xinput196 wb_rstn_i VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_12
Xinput197 wb_sel_i[0] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__clkbuf_1
Xinput198 wb_sel_i[1] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__clkbuf_1
Xinput199 wb_sel_i[2] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput2 debug_oeb VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
Xinput20 mask_rev_in[24] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput200 wb_sel_i[3] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput201 wb_stb_i VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__clkbuf_4
Xinput202 wb_we_i VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__clkbuf_2
Xinput21 mask_rev_in[25] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput22 mask_rev_in[26] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput23 mask_rev_in[27] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput24 mask_rev_in[28] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput25 mask_rev_in[29] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xinput26 mask_rev_in[2] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput27 mask_rev_in[30] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput28 mask_rev_in[31] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput29 mask_rev_in[3] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
Xinput3 debug_out VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
Xinput30 mask_rev_in[4] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
Xinput31 mask_rev_in[5] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xinput32 mask_rev_in[6] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput33 mask_rev_in[7] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput34 mask_rev_in[8] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_2
Xinput35 mask_rev_in[9] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput36 mgmt_gpio_in[0] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_8
Xinput37 mgmt_gpio_in[10] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput38 mgmt_gpio_in[11] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_6
Xinput39 mgmt_gpio_in[12] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput4 mask_rev_in[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xinput40 mgmt_gpio_in[13] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
Xinput41 mgmt_gpio_in[14] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput42 mgmt_gpio_in[15] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput43 mgmt_gpio_in[16] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput44 mgmt_gpio_in[17] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_1
Xinput45 mgmt_gpio_in[18] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
Xinput46 mgmt_gpio_in[19] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__clkbuf_1
Xinput47 mgmt_gpio_in[1] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_4
Xinput48 mgmt_gpio_in[20] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
Xinput49 mgmt_gpio_in[21] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_4
Xinput5 mask_rev_in[10] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
Xinput50 mgmt_gpio_in[22] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_4
Xinput51 mgmt_gpio_in[23] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_2
Xinput52 mgmt_gpio_in[24] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput53 mgmt_gpio_in[25] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_4
Xinput54 mgmt_gpio_in[26] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput55 mgmt_gpio_in[27] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput56 mgmt_gpio_in[28] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput57 mgmt_gpio_in[29] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput58 mgmt_gpio_in[2] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_12
Xinput59 mgmt_gpio_in[30] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
Xinput6 mask_rev_in[11] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
Xinput60 mgmt_gpio_in[31] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__clkbuf_1
Xinput61 mgmt_gpio_in[32] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_4
Xinput62 mgmt_gpio_in[33] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
Xinput63 mgmt_gpio_in[34] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_6
Xinput64 mgmt_gpio_in[35] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
Xinput65 mgmt_gpio_in[36] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
Xinput66 mgmt_gpio_in[37] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_4
Xinput67 mgmt_gpio_in[3] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_12
Xinput68 mgmt_gpio_in[5] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_4
Xinput69 mgmt_gpio_in[6] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_2
Xinput7 mask_rev_in[12] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
Xinput70 mgmt_gpio_in[7] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_1
Xinput71 mgmt_gpio_in[8] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__clkbuf_2
Xinput72 mgmt_gpio_in[9] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_1
Xinput73 pad_flash_io0_di VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__clkbuf_1
Xinput74 pad_flash_io1_di VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_2
Xinput75 porb VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_12
Xinput76 qspi_enabled VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_6
Xinput77 ser_tx VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_4
Xinput78 spi_csb VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_6
Xinput79 spi_enabled VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__buf_6
Xinput8 mask_rev_in[13] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
Xinput80 spi_sck VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__buf_6
Xinput81 spi_sdo VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__buf_6
Xinput82 spi_sdoenb VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_4
Xinput83 spimemio_flash_clk VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_6
Xinput84 spimemio_flash_csb VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_4
Xinput85 spimemio_flash_io0_do VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_4
Xinput86 spimemio_flash_io0_oeb VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_6
Xinput87 spimemio_flash_io1_do VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_6
Xinput88 spimemio_flash_io1_oeb VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_6
Xinput89 spimemio_flash_io2_do VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__clkbuf_4
Xinput9 mask_rev_in[14] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xinput90 spimemio_flash_io2_oeb VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_2
Xinput91 spimemio_flash_io3_do VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_4
Xinput92 spimemio_flash_io3_oeb VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__buf_2
Xinput93 sram_ro_data[0] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
Xinput94 sram_ro_data[10] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput95 sram_ro_data[11] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
Xinput96 sram_ro_data[12] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
Xinput97 sram_ro_data[13] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
Xinput98 sram_ro_data[14] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
Xinput99 sram_ro_data[15] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
Xnet299_2 clknet_2_3_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR net380 sky130_fd_sc_hd__inv_4
Xnet299_3 clknet_2_0_0_mgmt_gpio_in[4] VGND VGND VPWR VPWR net381 sky130_fd_sc_hd__inv_4
Xoutput203 net203 VGND VGND VPWR VPWR debug_in sky130_fd_sc_hd__buf_2
Xoutput204 net204 VGND VGND VPWR VPWR irq[0] sky130_fd_sc_hd__buf_2
Xoutput205 net205 VGND VGND VPWR VPWR irq[1] sky130_fd_sc_hd__buf_2
Xoutput206 net206 VGND VGND VPWR VPWR irq[2] sky130_fd_sc_hd__buf_2
Xoutput207 net207 VGND VGND VPWR VPWR mgmt_gpio_oeb[0] sky130_fd_sc_hd__buf_2
Xoutput208 net208 VGND VGND VPWR VPWR mgmt_gpio_oeb[10] sky130_fd_sc_hd__buf_2
Xoutput209 net209 VGND VGND VPWR VPWR mgmt_gpio_oeb[11] sky130_fd_sc_hd__buf_2
Xoutput210 net210 VGND VGND VPWR VPWR mgmt_gpio_oeb[12] sky130_fd_sc_hd__buf_2
Xoutput211 net211 VGND VGND VPWR VPWR mgmt_gpio_oeb[13] sky130_fd_sc_hd__buf_2
Xoutput212 net212 VGND VGND VPWR VPWR mgmt_gpio_oeb[14] sky130_fd_sc_hd__buf_2
Xoutput213 net213 VGND VGND VPWR VPWR mgmt_gpio_oeb[15] sky130_fd_sc_hd__buf_2
Xoutput214 net214 VGND VGND VPWR VPWR mgmt_gpio_oeb[16] sky130_fd_sc_hd__buf_2
Xoutput215 net215 VGND VGND VPWR VPWR mgmt_gpio_oeb[17] sky130_fd_sc_hd__buf_2
Xoutput216 net216 VGND VGND VPWR VPWR mgmt_gpio_oeb[18] sky130_fd_sc_hd__buf_2
Xoutput217 net217 VGND VGND VPWR VPWR mgmt_gpio_oeb[19] sky130_fd_sc_hd__buf_2
Xoutput218 net218 VGND VGND VPWR VPWR mgmt_gpio_oeb[1] sky130_fd_sc_hd__buf_2
Xoutput219 net219 VGND VGND VPWR VPWR mgmt_gpio_oeb[20] sky130_fd_sc_hd__buf_2
Xoutput220 net220 VGND VGND VPWR VPWR mgmt_gpio_oeb[21] sky130_fd_sc_hd__buf_2
Xoutput221 net221 VGND VGND VPWR VPWR mgmt_gpio_oeb[22] sky130_fd_sc_hd__buf_2
Xoutput222 net222 VGND VGND VPWR VPWR mgmt_gpio_oeb[23] sky130_fd_sc_hd__buf_2
Xoutput223 net223 VGND VGND VPWR VPWR mgmt_gpio_oeb[24] sky130_fd_sc_hd__buf_2
Xoutput224 net224 VGND VGND VPWR VPWR mgmt_gpio_oeb[25] sky130_fd_sc_hd__buf_2
Xoutput225 net225 VGND VGND VPWR VPWR mgmt_gpio_oeb[26] sky130_fd_sc_hd__buf_2
Xoutput226 net226 VGND VGND VPWR VPWR mgmt_gpio_oeb[27] sky130_fd_sc_hd__buf_2
Xoutput227 net227 VGND VGND VPWR VPWR mgmt_gpio_oeb[28] sky130_fd_sc_hd__buf_2
Xoutput228 net228 VGND VGND VPWR VPWR mgmt_gpio_oeb[29] sky130_fd_sc_hd__buf_2
Xoutput229 net229 VGND VGND VPWR VPWR mgmt_gpio_oeb[2] sky130_fd_sc_hd__buf_2
Xoutput230 net230 VGND VGND VPWR VPWR mgmt_gpio_oeb[30] sky130_fd_sc_hd__buf_2
Xoutput231 net231 VGND VGND VPWR VPWR mgmt_gpio_oeb[31] sky130_fd_sc_hd__buf_2
Xoutput232 net232 VGND VGND VPWR VPWR mgmt_gpio_oeb[32] sky130_fd_sc_hd__buf_2
Xoutput233 net233 VGND VGND VPWR VPWR mgmt_gpio_oeb[33] sky130_fd_sc_hd__buf_2
Xoutput234 net234 VGND VGND VPWR VPWR mgmt_gpio_oeb[34] sky130_fd_sc_hd__buf_2
Xoutput235 net235 VGND VGND VPWR VPWR mgmt_gpio_oeb[35] sky130_fd_sc_hd__buf_2
Xoutput236 net236 VGND VGND VPWR VPWR mgmt_gpio_oeb[36] sky130_fd_sc_hd__buf_2
Xoutput237 net237 VGND VGND VPWR VPWR mgmt_gpio_oeb[37] sky130_fd_sc_hd__buf_2
Xoutput238 net238 VGND VGND VPWR VPWR mgmt_gpio_oeb[3] sky130_fd_sc_hd__buf_2
Xoutput239 net239 VGND VGND VPWR VPWR mgmt_gpio_oeb[4] sky130_fd_sc_hd__buf_2
Xoutput240 net240 VGND VGND VPWR VPWR mgmt_gpio_oeb[5] sky130_fd_sc_hd__buf_2
Xoutput241 net241 VGND VGND VPWR VPWR mgmt_gpio_oeb[6] sky130_fd_sc_hd__buf_2
Xoutput242 net242 VGND VGND VPWR VPWR mgmt_gpio_oeb[7] sky130_fd_sc_hd__buf_2
Xoutput243 net243 VGND VGND VPWR VPWR mgmt_gpio_oeb[8] sky130_fd_sc_hd__buf_2
Xoutput244 net244 VGND VGND VPWR VPWR mgmt_gpio_oeb[9] sky130_fd_sc_hd__buf_2
Xoutput245 net245 VGND VGND VPWR VPWR mgmt_gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput246 net246 VGND VGND VPWR VPWR mgmt_gpio_out[1] sky130_fd_sc_hd__buf_2
Xoutput247 net247 VGND VGND VPWR VPWR mgmt_gpio_out[35] sky130_fd_sc_hd__buf_2
Xoutput248 net248 VGND VGND VPWR VPWR mgmt_gpio_out[36] sky130_fd_sc_hd__buf_2
Xoutput249 net249 VGND VGND VPWR VPWR mgmt_gpio_out[37] sky130_fd_sc_hd__buf_2
Xoutput250 net250 VGND VGND VPWR VPWR pad_flash_clk sky130_fd_sc_hd__clkbuf_1
Xoutput251 net251 VGND VGND VPWR VPWR pad_flash_clk_oeb sky130_fd_sc_hd__buf_2
Xoutput252 net252 VGND VGND VPWR VPWR pad_flash_csb sky130_fd_sc_hd__buf_2
Xoutput253 net253 VGND VGND VPWR VPWR pad_flash_csb_oeb sky130_fd_sc_hd__buf_2
Xoutput254 net254 VGND VGND VPWR VPWR pad_flash_io0_do sky130_fd_sc_hd__buf_2
Xoutput255 net255 VGND VGND VPWR VPWR pad_flash_io0_ieb sky130_fd_sc_hd__buf_2
Xoutput256 net256 VGND VGND VPWR VPWR pad_flash_io0_oeb sky130_fd_sc_hd__buf_2
Xoutput257 net257 VGND VGND VPWR VPWR pad_flash_io1_do sky130_fd_sc_hd__buf_2
Xoutput258 net258 VGND VGND VPWR VPWR pad_flash_io1_ieb sky130_fd_sc_hd__buf_2
Xoutput259 net259 VGND VGND VPWR VPWR pad_flash_io1_oeb sky130_fd_sc_hd__buf_2
Xoutput260 net260 VGND VGND VPWR VPWR pll90_sel[0] sky130_fd_sc_hd__buf_2
Xoutput261 net261 VGND VGND VPWR VPWR pll90_sel[1] sky130_fd_sc_hd__buf_2
Xoutput262 net262 VGND VGND VPWR VPWR pll90_sel[2] sky130_fd_sc_hd__buf_2
Xoutput263 net263 VGND VGND VPWR VPWR pll_bypass sky130_fd_sc_hd__buf_2
Xoutput264 net264 VGND VGND VPWR VPWR pll_dco_ena sky130_fd_sc_hd__buf_2
Xoutput265 net265 VGND VGND VPWR VPWR pll_div[0] sky130_fd_sc_hd__buf_2
Xoutput266 net266 VGND VGND VPWR VPWR pll_div[1] sky130_fd_sc_hd__buf_2
Xoutput267 net267 VGND VGND VPWR VPWR pll_div[2] sky130_fd_sc_hd__buf_2
Xoutput268 net268 VGND VGND VPWR VPWR pll_div[3] sky130_fd_sc_hd__buf_2
Xoutput269 net269 VGND VGND VPWR VPWR pll_div[4] sky130_fd_sc_hd__buf_2
Xoutput270 net270 VGND VGND VPWR VPWR pll_ena sky130_fd_sc_hd__buf_2
Xoutput271 net271 VGND VGND VPWR VPWR pll_sel[0] sky130_fd_sc_hd__buf_2
Xoutput272 net272 VGND VGND VPWR VPWR pll_sel[1] sky130_fd_sc_hd__buf_2
Xoutput273 net273 VGND VGND VPWR VPWR pll_sel[2] sky130_fd_sc_hd__buf_2
Xoutput274 net274 VGND VGND VPWR VPWR pll_trim[0] sky130_fd_sc_hd__buf_2
Xoutput275 net275 VGND VGND VPWR VPWR pll_trim[10] sky130_fd_sc_hd__buf_2
Xoutput276 net276 VGND VGND VPWR VPWR pll_trim[11] sky130_fd_sc_hd__buf_2
Xoutput277 net277 VGND VGND VPWR VPWR pll_trim[12] sky130_fd_sc_hd__buf_2
Xoutput278 net278 VGND VGND VPWR VPWR pll_trim[13] sky130_fd_sc_hd__buf_2
Xoutput279 net279 VGND VGND VPWR VPWR pll_trim[14] sky130_fd_sc_hd__buf_2
Xoutput280 net280 VGND VGND VPWR VPWR pll_trim[15] sky130_fd_sc_hd__buf_2
Xoutput281 net281 VGND VGND VPWR VPWR pll_trim[16] sky130_fd_sc_hd__buf_2
Xoutput282 net282 VGND VGND VPWR VPWR pll_trim[17] sky130_fd_sc_hd__buf_2
Xoutput283 net283 VGND VGND VPWR VPWR pll_trim[18] sky130_fd_sc_hd__buf_2
Xoutput284 net284 VGND VGND VPWR VPWR pll_trim[19] sky130_fd_sc_hd__buf_2
Xoutput285 net285 VGND VGND VPWR VPWR pll_trim[1] sky130_fd_sc_hd__buf_2
Xoutput286 net286 VGND VGND VPWR VPWR pll_trim[20] sky130_fd_sc_hd__buf_2
Xoutput287 net287 VGND VGND VPWR VPWR pll_trim[21] sky130_fd_sc_hd__buf_2
Xoutput288 net288 VGND VGND VPWR VPWR pll_trim[22] sky130_fd_sc_hd__buf_2
Xoutput289 net289 VGND VGND VPWR VPWR pll_trim[23] sky130_fd_sc_hd__buf_2
Xoutput290 net290 VGND VGND VPWR VPWR pll_trim[24] sky130_fd_sc_hd__buf_2
Xoutput291 net291 VGND VGND VPWR VPWR pll_trim[25] sky130_fd_sc_hd__buf_2
Xoutput292 net292 VGND VGND VPWR VPWR pll_trim[2] sky130_fd_sc_hd__buf_2
Xoutput293 net293 VGND VGND VPWR VPWR pll_trim[3] sky130_fd_sc_hd__buf_2
Xoutput294 net294 VGND VGND VPWR VPWR pll_trim[4] sky130_fd_sc_hd__buf_2
Xoutput295 net295 VGND VGND VPWR VPWR pll_trim[5] sky130_fd_sc_hd__buf_2
Xoutput296 net296 VGND VGND VPWR VPWR pll_trim[6] sky130_fd_sc_hd__buf_2
Xoutput297 net297 VGND VGND VPWR VPWR pll_trim[7] sky130_fd_sc_hd__buf_2
Xoutput298 net298 VGND VGND VPWR VPWR pll_trim[8] sky130_fd_sc_hd__buf_2
Xoutput299 net299 VGND VGND VPWR VPWR pll_trim[9] sky130_fd_sc_hd__buf_2
Xoutput300 net300 VGND VGND VPWR VPWR pwr_ctrl_out[0] sky130_fd_sc_hd__buf_2
Xoutput301 net301 VGND VGND VPWR VPWR pwr_ctrl_out[1] sky130_fd_sc_hd__buf_2
Xoutput302 net302 VGND VGND VPWR VPWR pwr_ctrl_out[2] sky130_fd_sc_hd__buf_2
Xoutput303 net303 VGND VGND VPWR VPWR pwr_ctrl_out[3] sky130_fd_sc_hd__buf_2
Xoutput304 net304 VGND VGND VPWR VPWR reset sky130_fd_sc_hd__buf_2
Xoutput305 net305 VGND VGND VPWR VPWR ser_rx sky130_fd_sc_hd__buf_2
Xoutput306 net306 VGND VGND VPWR VPWR serial_clock sky130_fd_sc_hd__clkbuf_1
Xoutput307 net307 VGND VGND VPWR VPWR serial_data_1 sky130_fd_sc_hd__buf_2
Xoutput308 net308 VGND VGND VPWR VPWR serial_data_2 sky130_fd_sc_hd__buf_2
Xoutput309 net309 VGND VGND VPWR VPWR serial_load sky130_fd_sc_hd__buf_2
Xoutput310 net310 VGND VGND VPWR VPWR serial_resetn sky130_fd_sc_hd__buf_2
Xoutput311 net311 VGND VGND VPWR VPWR spi_sdi sky130_fd_sc_hd__buf_2
Xoutput312 net312 VGND VGND VPWR VPWR spimemio_flash_io0_di sky130_fd_sc_hd__buf_2
Xoutput313 net313 VGND VGND VPWR VPWR spimemio_flash_io1_di sky130_fd_sc_hd__buf_2
Xoutput314 net314 VGND VGND VPWR VPWR spimemio_flash_io2_di sky130_fd_sc_hd__buf_2
Xoutput315 net315 VGND VGND VPWR VPWR spimemio_flash_io3_di sky130_fd_sc_hd__buf_2
Xoutput316 net316 VGND VGND VPWR VPWR sram_ro_addr[0] sky130_fd_sc_hd__buf_2
Xoutput317 net317 VGND VGND VPWR VPWR sram_ro_addr[1] sky130_fd_sc_hd__buf_2
Xoutput318 net318 VGND VGND VPWR VPWR sram_ro_addr[2] sky130_fd_sc_hd__buf_2
Xoutput319 net319 VGND VGND VPWR VPWR sram_ro_addr[3] sky130_fd_sc_hd__buf_2
Xoutput320 net320 VGND VGND VPWR VPWR sram_ro_addr[4] sky130_fd_sc_hd__buf_2
Xoutput321 net321 VGND VGND VPWR VPWR sram_ro_addr[5] sky130_fd_sc_hd__buf_2
Xoutput322 net322 VGND VGND VPWR VPWR sram_ro_addr[6] sky130_fd_sc_hd__buf_2
Xoutput323 net323 VGND VGND VPWR VPWR sram_ro_addr[7] sky130_fd_sc_hd__buf_2
Xoutput324 net324 VGND VGND VPWR VPWR sram_ro_clk sky130_fd_sc_hd__buf_2
Xoutput325 net325 VGND VGND VPWR VPWR sram_ro_csb sky130_fd_sc_hd__buf_2
Xoutput326 net326 VGND VGND VPWR VPWR wb_ack_o sky130_fd_sc_hd__buf_2
Xoutput327 net327 VGND VGND VPWR VPWR wb_dat_o[0] sky130_fd_sc_hd__buf_2
Xoutput328 net328 VGND VGND VPWR VPWR wb_dat_o[10] sky130_fd_sc_hd__buf_2
Xoutput329 net329 VGND VGND VPWR VPWR wb_dat_o[11] sky130_fd_sc_hd__buf_2
Xoutput330 net330 VGND VGND VPWR VPWR wb_dat_o[12] sky130_fd_sc_hd__buf_2
Xoutput331 net331 VGND VGND VPWR VPWR wb_dat_o[13] sky130_fd_sc_hd__buf_2
Xoutput332 net332 VGND VGND VPWR VPWR wb_dat_o[14] sky130_fd_sc_hd__buf_2
Xoutput333 net333 VGND VGND VPWR VPWR wb_dat_o[15] sky130_fd_sc_hd__buf_2
Xoutput334 net334 VGND VGND VPWR VPWR wb_dat_o[16] sky130_fd_sc_hd__buf_2
Xoutput335 net335 VGND VGND VPWR VPWR wb_dat_o[17] sky130_fd_sc_hd__buf_2
Xoutput336 net336 VGND VGND VPWR VPWR wb_dat_o[18] sky130_fd_sc_hd__buf_2
Xoutput337 net337 VGND VGND VPWR VPWR wb_dat_o[19] sky130_fd_sc_hd__buf_2
Xoutput338 net338 VGND VGND VPWR VPWR wb_dat_o[1] sky130_fd_sc_hd__buf_2
Xoutput339 net339 VGND VGND VPWR VPWR wb_dat_o[20] sky130_fd_sc_hd__buf_2
Xoutput340 net340 VGND VGND VPWR VPWR wb_dat_o[21] sky130_fd_sc_hd__buf_2
Xoutput341 net341 VGND VGND VPWR VPWR wb_dat_o[22] sky130_fd_sc_hd__buf_2
Xoutput342 net342 VGND VGND VPWR VPWR wb_dat_o[23] sky130_fd_sc_hd__buf_2
Xoutput343 net343 VGND VGND VPWR VPWR wb_dat_o[24] sky130_fd_sc_hd__buf_2
Xoutput344 net344 VGND VGND VPWR VPWR wb_dat_o[25] sky130_fd_sc_hd__buf_2
Xoutput345 net345 VGND VGND VPWR VPWR wb_dat_o[26] sky130_fd_sc_hd__buf_2
Xoutput346 net346 VGND VGND VPWR VPWR wb_dat_o[27] sky130_fd_sc_hd__buf_2
Xoutput347 net347 VGND VGND VPWR VPWR wb_dat_o[28] sky130_fd_sc_hd__buf_2
Xoutput348 net348 VGND VGND VPWR VPWR wb_dat_o[29] sky130_fd_sc_hd__buf_2
Xoutput349 net349 VGND VGND VPWR VPWR wb_dat_o[2] sky130_fd_sc_hd__buf_2
Xoutput350 net350 VGND VGND VPWR VPWR wb_dat_o[30] sky130_fd_sc_hd__buf_2
Xoutput351 net351 VGND VGND VPWR VPWR wb_dat_o[31] sky130_fd_sc_hd__buf_2
Xoutput352 net352 VGND VGND VPWR VPWR wb_dat_o[3] sky130_fd_sc_hd__buf_2
Xoutput353 net353 VGND VGND VPWR VPWR wb_dat_o[4] sky130_fd_sc_hd__buf_2
Xoutput354 net354 VGND VGND VPWR VPWR wb_dat_o[5] sky130_fd_sc_hd__buf_2
Xoutput355 net355 VGND VGND VPWR VPWR wb_dat_o[6] sky130_fd_sc_hd__buf_2
Xoutput356 net356 VGND VGND VPWR VPWR wb_dat_o[7] sky130_fd_sc_hd__buf_2
Xoutput357 net357 VGND VGND VPWR VPWR wb_dat_o[8] sky130_fd_sc_hd__buf_2
Xoutput358 net358 VGND VGND VPWR VPWR wb_dat_o[9] sky130_fd_sc_hd__buf_2
Xrepeater359 \cdata[4]\ VGND VGND VPWR VPWR net359 sky130_fd_sc_hd__buf_12
Xrepeater360 \cdata[4]\ VGND VGND VPWR VPWR net360 sky130_fd_sc_hd__buf_12
Xrepeater361 \cdata[3]\ VGND VGND VPWR VPWR net361 sky130_fd_sc_hd__buf_12
Xrepeater362 \cdata[3]\ VGND VGND VPWR VPWR net362 sky130_fd_sc_hd__buf_12
Xrepeater363 \cdata[2]\ VGND VGND VPWR VPWR net363 sky130_fd_sc_hd__buf_12
Xrepeater364 \cdata[2]\ VGND VGND VPWR VPWR net364 sky130_fd_sc_hd__buf_12
Xrepeater365 \cdata[1]\ VGND VGND VPWR VPWR net365 sky130_fd_sc_hd__buf_12
Xrepeater366 \cdata[1]\ VGND VGND VPWR VPWR net366 sky130_fd_sc_hd__buf_12
Xrepeater367 \cdata[0]\ VGND VGND VPWR VPWR net367 sky130_fd_sc_hd__buf_12
Xrepeater368 \cdata[0]\ VGND VGND VPWR VPWR net368 sky130_fd_sc_hd__buf_12
Xrepeater369 net370 VGND VGND VPWR VPWR net369 sky130_fd_sc_hd__buf_12
Xrepeater370 net75 VGND VGND VPWR VPWR net370 sky130_fd_sc_hd__buf_12
Xrepeater371 net373 VGND VGND VPWR VPWR net371 sky130_fd_sc_hd__buf_12
Xrepeater372 net373 VGND VGND VPWR VPWR net372 sky130_fd_sc_hd__buf_12
Xrepeater373 net374 VGND VGND VPWR VPWR net373 sky130_fd_sc_hd__buf_12
Xrepeater374 net375 VGND VGND VPWR VPWR net374 sky130_fd_sc_hd__buf_12
Xrepeater375 net75 VGND VGND VPWR VPWR net375 sky130_fd_sc_hd__buf_12
Xrepeater376 net377 VGND VGND VPWR VPWR net376 sky130_fd_sc_hd__buf_12
Xrepeater377 net75 VGND VGND VPWR VPWR net377 sky130_fd_sc_hd__buf_12

.ends
.end
