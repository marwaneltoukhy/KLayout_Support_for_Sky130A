* Extracted by KLayout on : 23/12/2021 16:56

.SUBCKT digital_pll osc clockp[0] clockp[1] div[0] VPWR div[1] div[2]
+ ext_trim[24] div[3] div[4] ext_trim[23] resetb enable dco ext_trim[0]
+ ext_trim[25] ext_trim[1] ext_trim[13] ext_trim[22] ext_trim[11] ext_trim[12]
+ ext_trim[14] ext_trim[2] ext_trim[21] ext_trim[18] ext_trim[10] ext_trim[9]
+ ext_trim[3] ext_trim[15] ext_trim[5] ext_trim[19] ext_trim[20] ext_trim[4]
+ ext_trim[6] ext_trim[17] ext_trim[16] ext_trim[7] ext_trim[8] VGND
X$1 VPWR osc VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2 VGND \$25 \$14 \$12 osc VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$3 VPWR VGND clockp[0] VPWR \$12 VGND sky130_fd_sc_hd__buf_2
X$4 VPWR VGND \$11 VPWR \$4 \$9 VGND sky130_fd_sc_hd__nor2_2
X$5 VPWR VPWR \$11 \$29 \$9 VGND \$4 VGND sky130_fd_sc_hd__a21oi_2
X$6 VGND \$96 \$9 \$11 \$49 \$4 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$7 VPWR \$18 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$8 VGND \$5 \$71 \$12 \$73 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9 VPWR VGND dco VPWR \$5 \$164 VGND sky130_fd_sc_hd__nor2_2
X$10 VPWR \$52 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$11 VPWR \$94 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$12 VPWR \$50 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$13 VPWR \$95 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$14 VPWR \$7 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$15 VPWR \$121 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$16 VPWR \$143 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$17 VPWR \$142 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$18 VPWR \$67 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$19 VPWR \$133 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$20 VPWR \$132 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$21 VPWR \$32 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$22 VPWR \$25 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$23 VPWR \$35 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$24 VPWR \$65 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$25 VPWR \$80 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$26 VPWR \$147 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$27 VPWR \$24 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$28 VPWR \$150 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$29 VPWR \$23 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$30 VPWR \$106 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$31 VGND clockp[1] \$169 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$32 VGND \$7 \$11 \$12 \$53 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$33 VGND \$37 \$63 \$64 \$31 \$8 VPWR VPWR VGND sky130_fd_sc_hd__and4_2
X$34 VGND \$24 \$8 \$12 \$16 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$35 VPWR \$16 VPWR VGND \$37 \$8 VGND sky130_fd_sc_hd__or2_2
X$36 VGND \$8 \$31 \$30 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$37 VGND \$11 \$9 \$19 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$38 VGND \$18 \$9 \$12 \$19 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$39 VPWR \$36 VPWR VGND \$20 \$10 \$21 VGND sky130_fd_sc_hd__or3_2
X$40 VPWR VGND VPWR \$10 \$15 VGND sky130_fd_sc_hd__inv_2
X$41 VGND \$27 \$15 \$45 \$21 \$10 \$13 VPWR VPWR VGND sky130_fd_sc_hd__o221a_2
X$42 VPWR \$10 VGND \$21 \$60 VPWR \$36 VGND sky130_fd_sc_hd__o21ai_2
X$43 VPWR VGND VPWR \$36 \$11 VGND sky130_fd_sc_hd__inv_2
X$44 VGND \$35 \$38 \$12 \$14 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$45 VGND \$12 \$139 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$46 VGND \$147 \$113 \$12 \$108 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$47 VGND \$143 \$144 \$12 \$137 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$48 VGND \$94 \$45 \$12 \$89 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$49 VGND \$23 \$15 \$12 \$22 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$50 VGND \$95 \$82 \$12 \$81 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$51 VGND \$80 \$77 \$12 \$104 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$52 VGND \$150 \$158 \$12 \$146 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$53 VGND \$65 \$42 \$12 \$38 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$54 VGND \$106 \$70 \$12 \$110 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$55 VGND \$50 \$34 \$12 \$51 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$56 VGND \$67 \$75 \$12 \$74 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$57 VGND \$142 \$166 \$12 \$165 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$58 VGND \$32 \$31 \$12 \$30 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$59 VGND \$52 \$63 \$12 \$56 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$60 VGND \$133 \$131 \$12 \$130 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$61 VGND \$121 \$126 \$12 \$115 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$62 VGND \$132 \$97 \$12 \$120 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$63 VPWR \$22 VPWR VGND \$13 \$62 VGND sky130_fd_sc_hd__or2_2
X$64 VGND \$41 \$34 \$15 \$34 \$15 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$65 VGND \$15 \$34 \$51 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$66 VGND \$46 \$15 \$44 \$41 \$34 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$67 VGND \$39 div[0] \$43 \$33 div[1] \$47 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$68 VPWR VGND VPWR \$59 div[0] VGND sky130_fd_sc_hd__inv_2
X$69 VPWR div[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$70 VPWR div[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$71 VPWR \$53 VPWR VGND \$60 \$20 \$27 \$62 VGND sky130_fd_sc_hd__a31o_2
X$72 VPWR VGND VPWR \$55 \$20 VGND sky130_fd_sc_hd__inv_2
X$73 VGND \$89 \$97 \$55 \$70 \$21 \$37 VPWR VPWR VGND sky130_fd_sc_hd__a311o_2
X$74 VPWR VPWR \$21 \$40 \$61 VGND \$46 VGND sky130_fd_sc_hd__a21oi_2
X$75 VPWR VGND VPWR \$21 \$45 VGND sky130_fd_sc_hd__inv_2
X$76 VPWR VGND \$21 VPWR \$46 \$61 VGND sky130_fd_sc_hd__nor2_2
X$77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$79 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$80 VPWR \$312 VPWR \$283 VGND \$317 VGND sky130_fd_sc_hd__einvp_2
X$81 VPWR \$288 VPWR \$287 VGND \$315 VGND sky130_fd_sc_hd__einvp_2
X$82 VPWR \$315 VGND VPWR \$289 VGND sky130_fd_sc_hd__clkbuf_1
X$83 VPWR VPWR VGND \$317 \$288 VGND sky130_fd_sc_hd__clkinv_1
X$84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$85 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$87 VPWR \$295 VPWR \$301 VGND \$318 VGND sky130_fd_sc_hd__einvp_2
X$88 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$89 VPWR \$316 VPWR \$310 VGND \$313 VGND sky130_fd_sc_hd__einvp_2
X$90 VPWR VPWR VGND \$318 \$316 VGND sky130_fd_sc_hd__clkinv_1
X$91 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$93 VPWR ext_trim[8] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$94 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$95 VPWR ext_trim[7] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$96 VGND \$311 ext_trim[7] \$220 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$97 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$99 VPWR \$314 VPWR \$311 VGND \$282 VGND sky130_fd_sc_hd__einvp_2
X$100 VPWR \$286 VPWR \$302 VGND \$303 VGND sky130_fd_sc_hd__einvp_2
X$101 VGND \$310 ext_trim[17] \$240 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$102 VPWR ext_trim[17] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$103 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$105 VGND \$287 ext_trim[16] \$276 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$106 VPWR \$309 VPWR \$306 VGND \$305 VGND sky130_fd_sc_hd__einvp_2
X$107 VPWR ext_trim[16] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$108 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$111 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$113 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$114 VPWR VGND VPWR \$43 \$40 VGND sky130_fd_sc_hd__inv_2
X$115 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$116 VGND \$48 \$44 \$29 \$44 VPWR \$29 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$118 VGND \$46 \$41 \$33 \$46 \$41 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2ai_2
X$119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$121 VPWR VGND VPWR \$37 \$27 VGND sky130_fd_sc_hd__inv_2
X$122 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$123 VGND \$27 \$38 \$42 \$38 VPWR \$42 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$124 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$127 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$128 VPWR VPWR \$39 \$33 VGND div[1] VGND sky130_fd_sc_hd__nand2_2
X$129 VGND \$57 \$54 \$58 \$47 \$40 \$59 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_2
X$130 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$131 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$132 VPWR VGND VPWR \$49 \$44 VGND sky130_fd_sc_hd__inv_2
X$133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$134 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$135 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$137 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$138 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$139 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$140 VGND \$63 \$31 \$56 \$27 \$37 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$141 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$143 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$145 VPWR div[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$147 VPWR \$69 VPWR \$66 VGND \$48 div[2] \$58 VGND sky130_fd_sc_hd__o211a_2
X$148 VPWR VPWR div[1] \$78 \$33 VGND \$47 VGND sky130_fd_sc_hd__a21oi_2
X$149 VGND \$70 \$71 \$73 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$151 VGND \$55 \$97 \$62 \$70 \$27 VPWR VPWR VGND sky130_fd_sc_hd__and4_2
X$152 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$155 VGND \$81 \$72 \$123 \$76 \$82 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$156 VPWR \$182 VPWR VGND \$79 \$77 \$82 VGND sky130_fd_sc_hd__or3_2
X$157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$159 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$162 VPWR div[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$163 VPWR div[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$164 VGND \$57 \$84 \$78 \$87 \$69 \$86 VPWR VPWR VGND sky130_fd_sc_hd__o221a_2
X$165 VPWR VGND VPWR \$84 \$58 VGND sky130_fd_sc_hd__inv_2
X$166 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$167 VPWR VGND \$70 VPWR \$88 \$71 VGND sky130_fd_sc_hd__nor2_2
X$168 VPWR VPWR VGND \$100 \$88 \$70 \$71 VGND sky130_fd_sc_hd__a21o_2
X$169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$171 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$172 VGND \$45 \$75 \$74 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$173 VPWR VGND VPWR \$61 \$75 VGND sky130_fd_sc_hd__inv_2
X$174 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$175 VGND \$64 \$101 \$79 \$54 \$91 \$92 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$176 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$177 VGND \$93 \$77 \$85 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$179 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$181 VPWR ext_trim[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$183 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$185 VPWR VPWR VGND \$216 \$238 VGND sky130_fd_sc_hd__clkbuf_2
X$186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$187 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$189 VPWR VPWR VGND \$213 \$218 VGND sky130_fd_sc_hd__clkinv_1
X$190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$191 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$192 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$193 VGND \$184 ext_trim[12] \$234 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$194 VGND \$290 \$214 \$158 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$196 VGND \$239 \$214 \$205 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$197 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$198 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$199 VGND \$219 ext_trim[14] \$235 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$201 VGND \$235 \$111 \$221 \$236 \$230 \$233 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$203 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$204 VGND \$240 \$233 \$221 \$111 \$131 \$236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$205 VPWR \$111 VPWR VGND \$241 \$205 \$221 VGND sky130_fd_sc_hd__or3_2
X$206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$207 VPWR ext_trim[21] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$208 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$209 VPWR VPWR VGND \$232 \$207 VGND sky130_fd_sc_hd__clkbuf_2
X$210 VGND \$243 ext_trim[22] \$233 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$211 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$214 VGND \$258 ext_trim[2] \$214 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$216 VGND \$238 \$248 \$245 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$217 VPWR \$259 VGND VPWR \$238 VGND sky130_fd_sc_hd__clkbuf_1
X$218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$219 VPWR VPWR VGND \$260 \$249 VGND sky130_fd_sc_hd__clkinv_1
X$220 VGND \$246 \$249 \$247 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$221 VGND \$234 \$126 \$221 \$158 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$223 VPWR \$250 VPWR VGND \$244 \$158 VGND sky130_fd_sc_hd__or2_2
X$224 VGND \$261 \$205 \$221 \$126 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$225 VGND \$226 ext_trim[10] \$251 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$226 VPWR \$251 VPWR VGND \$244 \$190 VGND sky130_fd_sc_hd__or2_2
X$227 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$228 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$229 VPWR ext_trim[14] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$230 VGND \$233 \$252 \$111 \$221 \$153 \$158 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$231 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$232 VGND \$254 \$158 \$153 \$187 \$126 \$204 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$233 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$235 VGND \$262 ext_trim[21] \$254 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$236 VPWR \$232 VPWR \$271 VGND \$255 VGND sky130_fd_sc_hd__einvp_2
X$237 VPWR \$256 VPWR \$243 VGND \$257 VGND sky130_fd_sc_hd__einvp_2
X$238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$241 VGND \$289 \$283 \$312 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$242 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$244 VGND \$289 \$288 \$287 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$245 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$246 VPWR VPWR VGND \$312 \$307 VGND sky130_fd_sc_hd__clkbuf_2
X$247 VPWR VPWR VGND \$273 \$289 VGND sky130_fd_sc_hd__clkbuf_2
X$248 VGND \$307 \$301 \$295 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$249 VPWR ext_trim[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$251 VGND \$301 ext_trim[4] \$290 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$252 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$253 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$254 VPWR VPWR VGND \$295 \$246 VGND sky130_fd_sc_hd__clkbuf_2
X$255 VGND \$307 \$316 \$310 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$256 VPWR ext_trim[6] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$257 VGND \$299 ext_trim[6] \$250 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$258 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$260 VGND \$269 \$299 \$300 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$261 VPWR \$313 VGND VPWR \$307 VGND sky130_fd_sc_hd__clkbuf_1
X$262 VGND \$306 ext_trim[8] \$261 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$263 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$264 VPWR VPWR VGND \$300 \$308 VGND sky130_fd_sc_hd__clkbuf_2
X$265 VPWR \$300 VPWR \$299 VGND \$291 VGND sky130_fd_sc_hd__einvp_2
X$266 VGND \$308 \$311 \$314 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$267 VPWR VPWR VGND \$291 \$284 VGND sky130_fd_sc_hd__clkinv_1
X$268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$269 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$270 VGND \$302 ext_trim[20] \$229 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$271 VGND \$308 \$286 \$302 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$272 VPWR \$303 VGND VPWR \$308 VGND sky130_fd_sc_hd__clkbuf_1
X$273 VPWR ext_trim[20] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$274 VGND \$281 ext_trim[19] \$267 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$275 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$276 VPWR \$293 VPWR \$262 VGND \$304 VGND sky130_fd_sc_hd__einvp_2
X$277 VPWR ext_trim[19] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$279 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$280 VGND \$294 \$293 \$262 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$281 VPWR VPWR VGND \$314 \$294 VGND sky130_fd_sc_hd__clkbuf_2
X$282 VGND \$294 \$306 \$309 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$283 VPWR \$304 VGND VPWR \$294 VGND sky130_fd_sc_hd__clkbuf_1
X$284 VPWR VPWR VGND \$305 \$293 VGND sky130_fd_sc_hd__clkinv_1
X$285 VPWR VPWR VGND \$309 \$268 VGND sky130_fd_sc_hd__clkbuf_2
X$286 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$287 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$292 VPWR ext_trim[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$293 VGND \$197 ext_trim[0] \$182 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$294 VGND \$202 \$197 \$183 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$295 VPWR \$183 VPWR \$197 VGND \$175 VGND sky130_fd_sc_hd__einvp_2
X$296 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$297 VPWR \$176 VPWR \$193 VGND \$192 VGND sky130_fd_sc_hd__einvp_2
X$298 VGND \$202 \$176 \$193 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$299 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$301 VPWR VPWR \$181 VGND \$164 \$198 VGND sky130_fd_sc_hd__einvp_1
X$302 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$303 VPWR \$199 VPWR VGND \$184 \$164 VGND sky130_fd_sc_hd__or2_2
X$304 VGND \$171 \$199 \$181 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$305 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$306 VPWR \$181 VPWR \$184 VGND \$194 VGND sky130_fd_sc_hd__einvp_2
X$307 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$308 VGND \$171 \$185 \$186 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$309 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$311 VPWR VPWR VGND \$194 \$185 VGND sky130_fd_sc_hd__clkinv_1
X$312 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$313 VPWR \$185 VPWR \$186 VGND \$177 VGND sky130_fd_sc_hd__einvp_2
X$314 VGND \$193 ext_trim[13] \$203 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$315 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$316 VPWR \$195 VGND \$101 \$155 VPWR \$178 VGND sky130_fd_sc_hd__o21ai_2
X$317 VPWR \$203 VPWR VGND \$158 \$166 \$144 \$126 VGND sky130_fd_sc_hd__a31o_2
X$318 VPWR VGND VPWR \$156 \$144 VGND sky130_fd_sc_hd__inv_2
X$319 VPWR \$187 VPWR VGND \$166 \$144 VGND sky130_fd_sc_hd__or2_2
X$320 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$321 VPWR VGND VPWR \$161 \$187 VGND sky130_fd_sc_hd__inv_2
X$322 VPWR VGND VPWR \$195 \$166 VGND sky130_fd_sc_hd__inv_2
X$323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$324 VGND \$186 ext_trim[25] \$188 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$325 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$326 VGND \$188 \$190 \$172 \$187 \$126 \$204 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$327 VPWR VGND \$190 VPWR \$170 \$172 VGND sky130_fd_sc_hd__nor2_2
X$328 VPWR \$182 VPWR VGND \$204 \$126 VGND sky130_fd_sc_hd__or2_2
X$329 VPWR ext_trim[25] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$330 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$331 VPWR VGND VPWR \$111 \$126 VGND sky130_fd_sc_hd__inv_2
X$332 VPWR VGND VPWR \$172 \$205 VGND sky130_fd_sc_hd__inv_2
X$333 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$334 VPWR \$171 VPWR \$206 VGND \$200 VGND sky130_fd_sc_hd__einvp_2
X$335 VPWR VPWR VGND \$200 \$191 VGND sky130_fd_sc_hd__clkinv_1
X$336 VPWR \$191 VPWR \$180 VGND \$179 VGND sky130_fd_sc_hd__einvp_2
X$337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$338 VGND \$174 \$206 \$171 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$339 VGND \$174 \$191 \$180 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$340 VPWR \$201 VPWR \$168 VGND \$196 VGND sky130_fd_sc_hd__einvp_2
X$341 VPWR \$196 VGND VPWR \$207 VGND sky130_fd_sc_hd__clkbuf_1
X$342 VPWR ext_trim[23] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$343 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$346 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$351 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$352 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$355 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$357 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$364 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$365 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$367 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$368 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$370 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$374 VGND \$283 ext_trim[3] \$244 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$375 VPWR ext_trim[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$376 VGND \$238 \$258 \$273 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$377 VPWR \$273 VPWR \$258 VGND \$277 VGND sky130_fd_sc_hd__einvp_2
X$378 VPWR \$248 VPWR \$245 VGND \$259 VGND sky130_fd_sc_hd__einvp_2
X$379 VPWR VPWR VGND \$277 \$248 VGND sky130_fd_sc_hd__clkinv_1
X$380 VPWR ext_trim[5] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$381 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$382 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$384 VGND \$265 ext_trim[5] \$278 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$385 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$386 VGND \$246 \$265 \$274 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$387 VPWR \$274 VPWR \$265 VGND \$260 VGND sky130_fd_sc_hd__einvp_2
X$388 VPWR \$249 VPWR \$247 VGND \$279 VGND sky130_fd_sc_hd__einvp_2
X$389 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$390 VGND \$278 \$126 \$221 \$190 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$391 VPWR \$279 VGND VPWR \$246 VGND sky130_fd_sc_hd__clkbuf_1
X$392 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$394 VPWR VGND VPWR \$214 \$244 \$221 \$126 VGND sky130_fd_sc_hd__o21a_2
X$395 VGND \$271 ext_trim[9] \$239 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$396 VPWR VPWR VGND \$274 \$269 VGND sky130_fd_sc_hd__clkbuf_2
X$397 VPWR ext_trim[10] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$398 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$399 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$400 VGND \$269 \$284 \$281 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$401 VPWR ext_trim[9] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$402 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$403 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$404 VPWR \$275 VGND VPWR \$269 VGND sky130_fd_sc_hd__clkbuf_1
X$405 VPWR VGND \$111 VPWR \$264 \$161 VGND sky130_fd_sc_hd__nor2_2
X$406 VPWR \$284 VPWR \$281 VGND \$275 VGND sky130_fd_sc_hd__einvp_2
X$407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$408 VGND \$247 ext_trim[18] \$264 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$409 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$410 VGND \$245 ext_trim[15] \$252 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$411 VPWR ext_trim[18] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$412 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$413 VPWR VPWR VGND \$282 \$286 VGND sky130_fd_sc_hd__clkinv_1
X$414 VGND \$252 \$111 \$187 \$236 \$241 \$254 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$415 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$416 VGND \$270 \$204 \$117 \$126 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$417 VPWR VPWR \$270 \$267 \$276 VGND VGND sky130_fd_sc_hd__and2_2
X$418 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$419 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$421 VPWR VPWR \$267 \$117 VGND \$111 VGND sky130_fd_sc_hd__nand2_2
X$422 VGND \$268 \$271 \$232 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$423 VPWR ext_trim[15] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$424 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$425 VPWR VPWR VGND \$255 \$256 VGND sky130_fd_sc_hd__clkinv_1
X$426 VGND \$268 \$256 \$243 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$427 VPWR \$257 VGND VPWR \$268 VGND sky130_fd_sc_hd__clkbuf_1
X$428 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$429 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$434 VPWR ext_trim[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$435 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$436 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$437 VPWR div[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$439 VPWR \$169 \$274 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$441 VPWR VPWR VGND \$175 \$176 VGND sky130_fd_sc_hd__clkinv_1
X$442 VPWR VGND VPWR \$114 \$113 VGND sky130_fd_sc_hd__inv_2
X$443 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$444 VPWR resetb VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$445 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$446 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$448 VPWR VPWR \$164 resetb VGND enable VGND sky130_fd_sc_hd__nand2_2
X$449 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$450 VPWR enable VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$451 VPWR \$139 \$181 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$456 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$457 VPWR \$177 VGND VPWR \$171 VGND sky130_fd_sc_hd__clkbuf_1
X$458 VPWR VGND VPWR \$160 \$155 VGND sky130_fd_sc_hd__inv_2
X$459 VPWR \$156 VGND \$76 \$137 VPWR \$167 VGND sky130_fd_sc_hd__o21ai_2
X$460 VPWR VGND VPWR \$152 \$151 VGND sky130_fd_sc_hd__inv_2
X$461 VGND \$151 \$152 \$167 \$123 \$160 \$155 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_2
X$462 VGND \$165 \$76 \$178 \$123 \$166 \$134 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$463 VGND \$151 \$144 \$101 \$102 \$156 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$464 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$465 VGND \$195 \$166 \$141 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$467 VGND \$124 \$141 \$151 \$140 \$161 \$101 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$468 VPWR \$178 VPWR VGND \$141 \$140 VGND sky130_fd_sc_hd__or2_2
X$469 VGND \$140 \$170 \$138 \$118 \$172 \$101 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$470 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$471 VGND \$153 \$131 \$138 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$472 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$473 VGND \$157 \$102 \$131 \$118 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$474 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$475 VPWR \$157 VPWR \$76 VGND \$101 \$153 \$149 VGND sky130_fd_sc_hd__o211a_2
X$476 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$478 VPWR VGND VPWR \$153 \$131 VGND sky130_fd_sc_hd__inv_2
X$479 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$480 VGND \$146 \$149 \$158 \$149 \$158 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2a_2
X$481 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$482 VPWR \$179 VGND VPWR \$174 VGND sky130_fd_sc_hd__clkbuf_1
X$483 VGND \$180 ext_trim[24] \$173 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$484 VGND \$168 ext_trim[23] \$159 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$485 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$486 VPWR \$159 VGND VPWR \$126 VGND sky130_fd_sc_hd__buf_1
X$487 VPWR ext_trim[24] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$492 VPWR div[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$493 VPWR div[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$494 VPWR VPWR \$57 \$119 VGND div[4] VGND sky130_fd_sc_hd__nand2_2
X$495 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$496 VGND \$112 \$91 div[4] \$119 \$122 \$114 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_2
X$497 VPWR \$112 VPWR VGND \$105 \$107 VGND sky130_fd_sc_hd__or2_2
X$498 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$499 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$500 VPWR VGND VPWR \$122 \$97 VGND sky130_fd_sc_hd__inv_2
X$501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$502 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$503 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$505 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$508 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$509 VPWR VGND VPWR \$123 \$76 VGND sky130_fd_sc_hd__inv_2
X$510 VPWR VGND VPWR \$127 \$124 VGND sky130_fd_sc_hd__inv_2
X$511 VGND \$128 \$111 \$101 \$102 \$126 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$512 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$513 VPWR VGND VPWR \$129 \$128 VGND sky130_fd_sc_hd__inv_2
X$514 VPWR VPWR \$134 \$141 VGND \$140 VGND sky130_fd_sc_hd__nand2_2
X$515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$516 VGND \$124 \$127 \$116 \$123 \$129 \$128 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_2
X$517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$518 VPWR VPWR \$135 \$138 VGND \$118 VGND sky130_fd_sc_hd__nand2_2
X$519 VGND \$130 \$76 \$145 \$123 \$131 \$135 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$520 VPWR \$145 VPWR VGND \$138 \$118 VGND sky130_fd_sc_hd__or2_2
X$521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$522 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$525 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$527 VGND \$48 div[2] \$69 div[3] \$99 VPWR VPWR VGND sky130_fd_sc_hd__a22oi_2
X$528 VPWR VGND VPWR \$87 \$66 VGND sky130_fd_sc_hd__inv_2
X$529 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$530 VGND \$99 \$100 \$96 \$100 VPWR \$96 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$531 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$533 VGND \$105 \$71 \$70 \$96 \$88 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$537 VPWR \$101 VPWR VGND \$91 \$86 VGND sky130_fd_sc_hd__or2_2
X$538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$539 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$541 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$542 VPWR VGND VPWR \$72 \$82 VGND sky130_fd_sc_hd__inv_2
X$543 VGND \$76 \$111 \$102 \$103 \$92 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$545 VGND \$123 \$104 \$98 \$76 \$93 VPWR VPWR VGND sky130_fd_sc_hd__o22ai_2
X$546 VGND \$98 \$72 \$85 \$72 VPWR \$85 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$548 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$551 VPWR \$66 VPWR VGND \$99 div[3] VGND sky130_fd_sc_hd__or2_2
X$552 VPWR VPWR VGND \$119 \$112 \$107 \$105 VGND sky130_fd_sc_hd__a21bo_2
X$553 VGND \$122 \$97 \$107 \$114 \$113 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$554 VGND \$97 \$113 \$108 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$555 VPWR VPWR \$122 \$120 \$109 VGND \$37 VGND sky130_fd_sc_hd__a21oi_2
X$556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$557 VGND \$27 \$97 \$109 \$55 \$70 \$110 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$558 VPWR VPWR \$109 \$55 VGND \$70 VGND sky130_fd_sc_hd__nand2_2
X$559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$560 VPWR VGND VPWR \$102 \$101 VGND sky130_fd_sc_hd__inv_2
X$561 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$562 VPWR \$111 VGND \$76 \$115 VPWR \$116 VGND sky130_fd_sc_hd__o21ai_2
X$563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$564 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$565 VPWR \$117 VPWR VGND \$103 \$93 \$72 VGND sky130_fd_sc_hd__or3_2
X$566 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$567 VGND \$118 \$72 \$85 \$101 \$93 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$569 VPWR VGND VPWR \$93 \$77 VGND sky130_fd_sc_hd__inv_2
X$570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$572 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$574 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$576 VGND \$223 ext_trim[1] \$212 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$577 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$578 VPWR \$216 VPWR \$223 VGND \$213 VGND sky130_fd_sc_hd__einvp_2
X$579 VPWR VPWR VGND \$183 \$224 VGND sky130_fd_sc_hd__clkbuf_2
X$580 VPWR \$192 VGND VPWR \$202 VGND sky130_fd_sc_hd__clkbuf_1
X$581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$582 VPWR \$218 VPWR \$219 VGND \$217 VGND sky130_fd_sc_hd__einvp_2
X$583 VPWR VPWR VGND \$181 \$202 VGND sky130_fd_sc_hd__clkbuf_2
X$584 VPWR VPWR VGND \$198 VGND sky130_fd_sc_hd__conb_1
X$585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$586 VGND \$212 \$156 \$166 \$126 \$214 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$588 VPWR \$220 VPWR VGND \$205 \$166 \$144 \$126 VGND sky130_fd_sc_hd__a31o_2
X$589 VPWR \$221 VPWR VGND \$195 \$144 VGND sky130_fd_sc_hd__or2_2
X$590 VPWR ext_trim[13] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$593 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$594 VPWR \$211 VPWR VGND \$117 \$156 \$195 VGND sky130_fd_sc_hd__or3_2
X$595 VPWR \$211 VPWR VGND \$153 \$236 VGND sky130_fd_sc_hd__or2_2
X$596 VPWR VGND VPWR \$190 \$211 VGND sky130_fd_sc_hd__inv_2
X$597 VPWR \$126 \$187 \$221 VGND VPWR \$173 VGND sky130_fd_sc_hd__and3_2
X$598 VPWR \$205 VPWR VGND \$131 \$158 VGND sky130_fd_sc_hd__or2_2
X$599 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$600 VPWR VPWR VGND \$215 \$174 VGND sky130_fd_sc_hd__clkbuf_2
X$601 VPWR \$215 VPWR \$226 VGND \$222 VGND sky130_fd_sc_hd__einvp_2
X$602 VGND \$207 \$201 \$168 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$605 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$606 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$607 VGND \$224 \$223 \$216 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$608 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$609 VGND \$224 \$218 \$219 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$610 VPWR \$217 VGND VPWR \$224 VGND sky130_fd_sc_hd__clkbuf_1
X$611 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$612 VGND \$206 ext_trim[11] \$225 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$613 VPWR ext_trim[11] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$614 VPWR ext_trim[12] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$617 VGND \$225 \$214 \$190 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$619 VPWR \$244 VPWR VGND \$187 \$126 VGND sky130_fd_sc_hd__or2_2
X$620 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$621 VPWR \$205 \$166 VGND \$156 VPWR \$230 \$111 VGND sky130_fd_sc_hd__or4_2
X$622 VGND \$229 \$156 \$166 \$158 \$173 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$624 VPWR \$204 VPWR VGND \$187 \$205 VGND sky130_fd_sc_hd__or2_2
X$625 VPWR VGND VPWR \$236 \$158 VGND sky130_fd_sc_hd__inv_2
X$626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$628 VGND \$207 \$226 \$215 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$629 VPWR VPWR VGND \$222 \$201 VGND sky130_fd_sc_hd__clkinv_1
X$630 VPWR ext_trim[22] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
.ENDS digital_pll

.SUBCKT sky130_fd_sc_hd__o22a_2 VGND X B1 B2 A2 A1 VPB VPWR VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=390000000000P PS=1270000U PD=1780000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=390000000000P AD=105000000000P PS=1780000U PD=1210000U
M$4 \$12 B2 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=235000000000P PS=1210000U PD=1470000U
M$5 \$4 A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=235000000000P AD=105000000000P PS=1470000U PD=1210000U
M$6 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=280000000000P PS=1210000U PD=2560000U
M$7 \$6 B1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$8 \$4 B2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=123500000000P PS=920000U PD=1030000U
M$9 \$6 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=87750000000P PS=1030000U PD=920000U
M$10 VGND A1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$11 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$12 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22a_2

.SUBCKT sky130_fd_sc_hd__o22ai_2 VGND B1 Y B2 A2 A1 VPWR VPB VNB
M$1 \$11 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 Y A2 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$11 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 VPWR A1 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=280000000000P PS=1270000U PD=2560000U
M$5 \$9 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$6 VPWR B1 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$9 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Y B2 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=280000000000P PS=1270000U PD=2560000U
M$9 \$3 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=182000000000P
+ AD=87750000000P PS=1860000U PD=920000U
M$10 Y B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 \$3 B2 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$12 Y B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=269750000000P PS=920000U PD=1480000U
M$13 \$3 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=269750000000P AD=87750000000P PS=1480000U PD=920000U
M$14 VGND A2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$3 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$16 VGND A1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o22ai_2

.SUBCKT sky130_fd_sc_hd__and4_2 VGND B C X A D VPWR VPB VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=74550000000P PS=1360000U PD=775000U
M$2 \$3 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74550000000P AD=77700000000P PS=775000U PD=790000U
M$3 VPWR C \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=77700000000P AD=58800000000P PS=790000U PD=700000U
M$4 VPWR D \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=279950000000P AD=58800000000P PS=1615000U PD=700000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=279950000000P AD=165000000000P PS=1615000U PD=1330000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=300000000000P PS=1330000U PD=2600000U
M$7 \$3 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=61950000000P PS=1360000U PD=715000U
M$8 \$9 B \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=61950000000P
+ AD=79800000000P PS=715000U PD=800000U
M$9 \$10 C \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=79800000000P
+ AD=69300000000P PS=800000U PD=750000U
M$10 \$11 D VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=175150000000P PS=750000U PD=1265000U
M$11 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=175150000000P AD=107250000000P PS=1265000U PD=980000U
M$12 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=195000000000P PS=980000U PD=1900000U
.ENDS sky130_fd_sc_hd__and4_2

.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 VGND A1_N A2_N Y B1 B2 VPWR VPB VNB
M$1 VPWR A1_N \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 \$6 A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A2_N \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$6 A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=400000000000P PS=1270000U PD=1800000U
M$5 VPWR \$6 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=400000000000P AD=135000000000P PS=1800000U PD=1270000U
M$6 Y \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=152500000000P PS=1270000U PD=1305000U
M$7 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=152500000000P AD=135000000000P PS=1305000U PD=1270000U
M$8 \$12 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 Y B2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 \$12 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$11 \$7 \$6 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=175500000000P
+ AD=87750000000P PS=1840000U PD=920000U
M$12 Y \$6 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=99125000000P PS=920000U PD=955000U
M$13 \$7 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=99125000000P AD=87750000000P PS=955000U PD=920000U
M$14 VGND B2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$7 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$16 VGND B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$17 VGND A1_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=182000000000P AD=87750000000P PS=1860000U PD=920000U
M$18 \$4 A2_N \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$19 \$6 A2_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$20 \$4 A1_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o2bb2ai_2

.SUBCKT sky130_fd_sc_hd__o211a_2 VPB C1 VPWR B1 VGND A2 A1 X VNB
M$1 \$3 C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 VPWR B1 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=367500000000P PS=1280000U PD=1735000U
M$3 \$3 A2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=367500000000P AD=105000000000P PS=1735000U PD=1210000U
M$4 \$12 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=195000000000P PS=1210000U PD=1390000U
M$5 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=140000000000P PS=1390000U PD=1280000U
M$6 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$7 VGND A2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=165350000000P AD=91000000000P PS=1820000U PD=930000U
M$8 \$7 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=104000000000P PS=930000U PD=970000U
M$9 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=104000000000P
+ AD=91000000000P PS=970000U PD=930000U
M$10 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=230750000000P PS=930000U PD=2010000U
M$11 \$3 C1 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=68250000000P PS=1830000U PD=860000U
M$12 \$13 B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=165350000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o211a_2

.SUBCKT sky130_fd_sc_hd__o2111ai_2 VGND D1 Y C1 B1 A2 A1 VPWR VPB VNB
M$1 \$13 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=295000000000P AD=140000000000P PS=2590000U PD=1280000U
M$2 Y A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$4 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=330000000000P PS=1280000U PD=2660000U
M$5 VPWR D1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$6 Y D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$7 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$8 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$9 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$10 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$11 \$9 B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=175500000000P AD=91000000000P PS=1840000U PD=930000U
M$12 \$7 B1 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$13 \$9 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$14 VGND A2 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$15 \$9 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=91000000000P PS=930000U PD=930000U
M$16 VGND A1 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=91000000000P AD=214500000000P PS=930000U PD=1960000U
M$17 \$4 D1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=224250000000P
+ AD=91000000000P PS=1990000U PD=930000U
M$18 Y D1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$19 \$4 C1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$20 \$7 C1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=191750000000P PS=930000U PD=1890000U
.ENDS sky130_fd_sc_hd__o2111ai_2

.SUBCKT sky130_fd_sc_hd__buf_2 VPB VGND X VPWR A VNB
M$1 VPWR A \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=149000000000P AD=166400000000P PS=1325000U PD=1800000U
M$2 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=149000000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=265000000000P PS=1270000U PD=2530000U
M$4 \$4 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=97000000000P PS=1360000U PD=975000U
M$5 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$6 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=172250000000P PS=920000U PD=1830000U
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__o221ai_2 VGND C1 Y B1 B2 A1 A2 VPWR VPB VNB
M$1 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=395000000000P PS=1270000U PD=1790000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=395000000000P AD=135000000000P PS=1790000U PD=1270000U
M$4 \$12 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 Y B2 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 \$12 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=175000000000P PS=1270000U PD=1350000U
M$7 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=135000000000P PS=1350000U PD=1270000U
M$8 \$13 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 Y A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$11 \$6 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$12 \$3 B2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$13 \$6 B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$14 \$3 B1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=113750000000P PS=920000U PD=1000000U
M$15 \$6 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=87750000000P PS=1000000U PD=920000U
M$16 VGND A2 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$17 \$6 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$18 VGND A1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$19 \$3 C1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$20 Y C1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221ai_2

.SUBCKT sky130_fd_sc_hd__a21bo_2 VPB VPWR VGND X B1_N A1 A2 VNB
M$1 \$9 \$8 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 \$3 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A2 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$4 VPWR B1_N \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=181500000000P AD=109200000000P PS=1510000U PD=1360000U
M$5 VPWR \$9 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=140000000000P PS=2520000U PD=1280000U
M$6 X \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=181500000000P PS=1280000U PD=1510000U
M$7 VGND \$8 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$8 \$9 A1 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=68250000000P PS=980000U PD=860000U
M$9 \$12 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=169000000000P PS=860000U PD=1820000U
M$10 VGND \$9 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=91000000000P PS=1820000U PD=930000U
M$11 X \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=108375000000P PS=930000U PD=1010000U
M$12 VGND B1_N \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=108375000000P AD=109200000000P PS=1010000U PD=1360000U
.ENDS sky130_fd_sc_hd__a21bo_2

.SUBCKT sky130_fd_sc_hd__a2bb2o_2 VGND X A1_N A2_N B1 VPWR B2 VPB VNB
M$1 \$6 \$4 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=97600000000P PS=1800000U PD=945000U
M$2 \$12 B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=97600000000P AD=86400000000P PS=945000U PD=910000U
M$3 VPWR B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$4 VPWR A1_N \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=186000000000P AD=67200000000P PS=1435000U PD=850000U
M$5 \$13 A2_N \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=67200000000P AD=169600000000P PS=850000U PD=1810000U
M$6 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=135000000000P PS=2530000U PD=1270000U
M$7 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=186000000000P PS=1270000U PD=1435000U
M$8 VGND A1_N \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=120100000000P AD=56700000000P PS=1085000U PD=690000U
M$9 \$4 A2_N VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=141750000000P PS=690000U PD=1095000U
M$10 VGND \$4 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=141750000000P AD=56700000000P PS=1095000U PD=690000U
M$11 \$6 B2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$12 \$5 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$13 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=87750000000P PS=1830000U PD=920000U
M$14 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=120100000000P PS=920000U PD=1085000U
.ENDS sky130_fd_sc_hd__a2bb2o_2

.SUBCKT sky130_fd_sc_hd__a22oi_2 VGND B2 B1 Y A1 A2 VPWR VPB VNB
M$1 \$10 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 VPWR A1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$10 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 VPWR A2 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 Y B2 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$10 B2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 Y B1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 \$10 B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$9 \$7 A1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$10 Y A1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 \$7 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$12 VGND A2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
M$13 \$3 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$14 VGND B2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$15 \$3 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$16 Y B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22oi_2

.SUBCKT sky130_fd_sc_hd__a311o_2 VGND X A3 A2 A1 B1 C1 VPWR VPB VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=240000000000P PS=1270000U PD=1480000U
M$3 VPWR A3 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=240000000000P AD=170000000000P PS=1480000U PD=1340000U
M$4 \$13 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=170000000000P AD=185000000000P PS=1340000U PD=1370000U
M$5 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=185000000000P AD=210000000000P PS=1370000U PD=1420000U
M$6 \$13 B1 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=210000000000P PS=1420000U PD=1420000U
M$7 \$15 C1 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=260000000000P PS=1420000U PD=2520000U
M$8 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=156000000000P PS=920000U PD=1130000U
M$10 VGND A3 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=156000000000P AD=110500000000P PS=1130000U PD=990000U
M$11 \$6 A2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=110500000000P AD=120250000000P PS=990000U PD=1020000U
M$12 \$5 A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=120250000000P AD=133250000000P PS=1020000U PD=1060000U
M$13 \$4 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=133250000000P AD=139750000000P PS=1060000U PD=1080000U
M$14 VGND C1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=169000000000P PS=1080000U PD=1820000U
.ENDS sky130_fd_sc_hd__a311o_2

.SUBCKT sky130_fd_sc_hd__a21oi_2 VPB VPWR A1 Y A2 VGND B1 VNB
M$1 \$5 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=140000000000P PS=2560000U PD=1280000U
M$2 VPWR A1 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 \$5 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=135000000000P PS=1280000U PD=1270000U
M$4 VPWR A2 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 \$5 B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Y B1 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=360000000000P PS=1270000U PD=2720000U
M$7 VGND A2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=185250000000P AD=89375000000P PS=1870000U PD=925000U
M$8 \$10 A1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=89375000000P
+ AD=91000000000P PS=925000U PD=930000U
M$9 Y A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=68250000000P PS=930000U PD=860000U
M$10 \$11 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=107250000000P PS=860000U PD=980000U
M$11 VGND B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=107250000000P
+ AD=87750000000P PS=980000U PD=920000U
M$12 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=260000000000P PS=920000U PD=2100000U
.ENDS sky130_fd_sc_hd__a21oi_2

.SUBCKT sky130_fd_sc_hd__a21o_2 VPB VPWR VGND X B1 A1 A2 VNB
M$1 \$7 B1 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$3 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=157500000000P PS=1280000U PD=1315000U
M$3 VPWR A2 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=260000000000P PS=1315000U PD=2520000U
M$4 VPWR \$7 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$5 X \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$6 VGND \$7 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=172250000000P
+ AD=91000000000P PS=1830000U PD=930000U
M$7 X \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=110500000000P PS=930000U PD=990000U
M$8 VGND B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=110500000000P AD=162500000000P PS=990000U PD=1150000U
M$9 \$7 A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=162500000000P AD=123500000000P PS=1150000U PD=1030000U
M$10 \$11 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=172250000000P PS=1030000U PD=1830000U
.ENDS sky130_fd_sc_hd__a21o_2

.SUBCKT sky130_fd_sc_hd__o221a_2 VGND C1 B1 B2 A2 A1 X VPB VPWR VNB
M$1 \$4 C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=325000000000P AD=165000000000P PS=2650000U PD=1330000U
M$2 VPWR B1 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=112500000000P PS=1330000U PD=1225000U
M$3 \$14 B2 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=112500000000P AD=387500000000P PS=1225000U PD=1775000U
M$4 \$4 A2 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=387500000000P AD=105000000000P PS=1775000U PD=1210000U
M$5 \$15 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=105000000000P AD=165000000000P PS=1210000U PD=1330000U
M$6 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=135000000000P PS=1330000U PD=1270000U
M$7 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 VGND A2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$9 \$7 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$10 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$11 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$12 \$4 C1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=237250000000P AD=87750000000P PS=2030000U PD=920000U
M$13 \$5 B1 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$14 \$7 B2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o221a_2

.SUBCKT sky130_fd_sc_hd__conb_1 VPB VPWR VGND HI VNB
R$1 VGND LO 0 sky130_fd_pr__res_generic_po
R$2 HI VPWR 0 sky130_fd_pr__res_generic_po
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__einvp_1 VPB VPWR Z VGND TE A VNB
M$1 VPWR TE \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=320750000000P AD=109200000000P PS=1685000U PD=1360000U
M$2 VPWR \$7 \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=320750000000P AD=182500000000P PS=1685000U PD=1365000U
M$3 \$9 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=182500000000P AD=270000000000P PS=1365000U PD=2540000U
M$4 \$7 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$5 VGND TE \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=97000000000P AD=235625000000P PS=975000U PD=1375000U
M$6 \$10 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=235625000000P
+ AD=175500000000P PS=1375000U PD=1840000U
.ENDS sky130_fd_sc_hd__einvp_1

.SUBCKT sky130_fd_sc_hd__o21a_2 VPB VGND VPWR X B1 A2 A1 VNB
M$1 VPWR \$6 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=137500000000P PS=2520000U PD=1275000U
M$2 X \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=400000000000P PS=1275000U PD=1800000U
M$3 VPWR B1 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=400000000000P AD=140000000000P PS=1800000U PD=1280000U
M$4 \$6 A2 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=160000000000P PS=1280000U PD=1320000U
M$5 \$11 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160000000000P AD=265000000000P PS=1320000U PD=2530000U
M$6 \$6 B1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=172250000000P
+ AD=91000000000P PS=1830000U PD=930000U
M$7 \$8 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=104000000000P PS=930000U PD=970000U
M$8 VGND A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=104000000000P AD=172250000000P PS=970000U PD=1830000U
M$9 VGND \$6 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=89375000000P PS=1820000U PD=925000U
M$10 X \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=89375000000P
+ AD=172250000000P PS=925000U PD=1830000U
.ENDS sky130_fd_sc_hd__o21a_2

.SUBCKT sky130_fd_sc_hd__or3_2 VPB C VPWR VGND X A B VNB
M$1 \$8 C \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$2 \$11 B \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$3 \$10 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=148250000000P PS=750000U PD=1340000U
M$4 VPWR \$8 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=148250000000P AD=135000000000P PS=1340000U PD=1270000U
M$5 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=315000000000P PS=1270000U PD=2630000U
M$6 \$8 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$7 VGND B \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$8 VGND A \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=101875000000P
+ AD=56700000000P PS=990000U PD=690000U
M$9 VGND \$8 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=101875000000P
+ AD=87750000000P PS=990000U PD=920000U
M$10 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=185250000000P PS=920000U PD=1870000U
.ENDS sky130_fd_sc_hd__or3_2

.SUBCKT sky130_fd_sc_hd__decap_8 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=2890000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=2890000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__or4_2 VPB C B VGND A VPWR X D VNB
M$1 \$5 D \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=69300000000P PS=1360000U PD=750000U
M$2 \$13 C \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=44100000000P PS=750000U PD=630000U
M$3 \$12 B \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$4 \$11 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=148250000000P PS=750000U PD=1340000U
M$5 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=148250000000P AD=135000000000P PS=1340000U PD=1270000U
M$6 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=2610000U
M$7 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=69300000000P PS=1360000U PD=750000U
M$8 \$5 C VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=56700000000P PS=750000U PD=690000U
M$9 VGND B \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=56700000000P PS=690000U PD=690000U
M$10 VGND A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=101875000000P AD=56700000000P PS=990000U PD=690000U
M$11 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=101875000000P AD=87750000000P PS=990000U PD=920000U
M$12 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=198250000000P PS=920000U PD=1910000U
.ENDS sky130_fd_sc_hd__or4_2

.SUBCKT sky130_fd_sc_hd__clkbuf_2 VPB VPWR VGND A X VNB
M$1 \$5 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=162500000000P PS=2530000U PD=1325000U
M$2 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=162500000000P AD=135000000000P PS=1325000U PD=1270000U
M$3 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$4 \$5 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=68250000000P PS=1370000U PD=745000U
M$5 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=68250000000P
+ AD=56700000000P PS=745000U PD=690000U
M$6 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__nand2_2 VPB VPWR Y B VGND A VNB
M$1 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$4 B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$6 VGND B \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$7 \$4 A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$8 Y A \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__and2_2 VPB VPWR A B X VGND VNB
M$1 VPWR A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=117600000000P AD=56700000000P PS=1400000U PD=690000U
M$2 VPWR B \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=166550000000P AD=56700000000P PS=1390000U PD=690000U
M$3 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=166550000000P AD=195000000000P PS=1390000U PD=1390000U
M$4 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=380000000000P PS=1390000U PD=2760000U
M$5 \$3 A \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=117600000000P
+ AD=56700000000P PS=1400000U PD=690000U
M$6 VGND B \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111800000000P
+ AD=56700000000P PS=1040000U PD=690000U
M$7 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=111800000000P
+ AD=126750000000P PS=1040000U PD=1040000U
M$8 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=126750000000P
+ AD=247000000000P PS=1040000U PD=2060000U
.ENDS sky130_fd_sc_hd__and2_2

.SUBCKT sky130_fd_sc_hd__einvp_2 VPB Z VPWR TE VGND A VNB
M$1 \$3 \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=244400000000P AD=126900000000P PS=2400000U PD=1210000U
M$2 \$3 \$6 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=160250000000P AD=126900000000P PS=1325000U PD=1210000U
M$3 \$3 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160250000000P AD=135000000000P PS=1325000U PD=1270000U
M$4 Z A \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$6 TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=166400000000P PS=1800000U PD=1800000U
M$6 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$7 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$8 \$6 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=97000000000P PS=1360000U PD=975000U
M$9 VGND TE \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=97000000000P
+ AD=87750000000P PS=975000U PD=920000U
M$10 \$5 TE VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__einvp_2

.SUBCKT sky130_fd_sc_hd__o311a_2 VGND X A1 A2 A3 B1 C1 VPWR VPB VNB
M$1 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=320000000000P AD=135000000000P PS=2640000U PD=1270000U
M$2 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=312500000000P PS=1270000U PD=1625000U
M$3 VPWR A1 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=312500000000P AD=175000000000P PS=1625000U PD=1350000U
M$4 \$14 A2 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=210000000000P PS=1350000U PD=1420000U
M$5 \$15 A3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=210000000000P AD=137500000000P PS=1420000U PD=1275000U
M$6 \$5 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=150000000000P PS=1275000U PD=1300000U
M$7 VPWR C1 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=150000000000P AD=260000000000P PS=1300000U PD=2520000U
M$8 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=208000000000P
+ AD=87750000000P PS=1940000U PD=920000U
M$9 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=203125000000P PS=920000U PD=1275000U
M$10 VGND A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=203125000000P AD=113750000000P PS=1275000U PD=1000000U
M$11 \$4 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=136500000000P PS=1000000U PD=1070000U
M$12 VGND A3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=136500000000P AD=118625000000P PS=1070000U PD=1015000U
M$13 \$4 B1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=118625000000P AD=68250000000P PS=1015000U PD=860000U
M$14 \$11 C1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=68250000000P AD=169000000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__o311a_2

.SUBCKT sky130_fd_sc_hd__and3_2 VPB A B C VGND VPWR X VNB
M$1 \$5 C VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74375000000P AD=150750000000P PS=815000U PD=1345000U
M$2 \$5 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$3 \$5 B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=74375000000P AD=56700000000P PS=815000U PD=690000U
M$4 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=150750000000P AD=135000000000P PS=1345000U PD=1270000U
M$5 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 \$5 A \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=44100000000P PS=1360000U PD=630000U
M$7 \$11 B \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=44100000000P
+ AD=53550000000P PS=630000U PD=675000U
M$8 VGND C \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=130400000000P AD=53550000000P PS=1105000U PD=675000U
M$9 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=130400000000P
+ AD=87750000000P PS=1105000U PD=920000U
M$10 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=178750000000P PS=920000U PD=1850000U
.ENDS sky130_fd_sc_hd__and3_2

.SUBCKT sky130_fd_sc_hd__einvn_4 VGND A Z TE_B VPWR VPB VNB
M$1 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 \$4 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=160250000000P PS=2520000U PD=1325000U
M$6 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=160250000000P AD=126900000000P PS=1325000U PD=1210000U
M$7 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$8 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$9 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=244400000000P PS=1210000U PD=2400000U
M$10 \$5 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$11 VGND \$4 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$12 \$5 \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$13 VGND \$4 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=105625000000P PS=920000U PD=975000U
M$14 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=105625000000P
+ AD=87750000000P PS=975000U PD=920000U
M$15 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$16 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$17 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=182000000000P PS=920000U PD=1860000U
M$18 \$4 TE_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=169000000000P PS=1820000U PD=1820000U
.ENDS sky130_fd_sc_hd__einvn_4

.SUBCKT sky130_fd_sc_hd__einvn_8 VGND A TE_B Z VPWR VPB VNB
M$1 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$8 A Z VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Z A \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$9 \$6 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=160250000000P PS=2520000U PD=1325000U
M$10 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=160250000000P AD=126900000000P PS=1325000U PD=1210000U
M$11 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$12 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$13 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$14 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$15 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$16 VPWR TE_B \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=126900000000P PS=1210000U PD=1210000U
M$17 \$8 TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=940000U
+ AS=126900000000P AD=244400000000P PS=1210000U PD=2400000U
M$18 \$6 TE_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=169000000000P PS=1820000U PD=1820000U
M$19 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$20 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$21 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$22 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$23 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$24 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$25 \$5 \$6 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$26 VGND \$6 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=105625000000P PS=920000U PD=975000U
M$27 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=105625000000P
+ AD=87750000000P PS=975000U PD=920000U
M$28 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$29 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$30 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$31 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$32 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$33 \$5 A Z VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$34 Z A \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=182000000000P PS=920000U PD=1860000U
.ENDS sky130_fd_sc_hd__einvn_8

.SUBCKT sky130_fd_sc_hd__o31a_2 VGND X A1 A2 A3 B1 VPWR VPB VNB
M$1 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=405000000000P AD=175000000000P PS=2810000U PD=1350000U
M$2 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=195000000000P PS=1350000U PD=1390000U
M$3 VPWR A1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=195000000000P AD=135000000000P PS=1390000U PD=1270000U
M$4 \$12 A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=165000000000P PS=1270000U PD=1330000U
M$5 \$13 A3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=212500000000P PS=1330000U PD=1425000U
M$6 \$5 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=212500000000P AD=340000000000P PS=1425000U PD=2680000U
M$7 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=263250000000P
+ AD=113750000000P PS=2110000U PD=1000000U
M$8 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=113750000000P
+ AD=126750000000P PS=1000000U PD=1040000U
M$9 VGND A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=87750000000P PS=1040000U PD=920000U
M$10 \$4 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=107250000000P PS=920000U PD=980000U
M$11 VGND A3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=107250000000P PS=980000U PD=980000U
M$12 \$4 B1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=201500000000P PS=980000U PD=1920000U
.ENDS sky130_fd_sc_hd__o31a_2

.SUBCKT sky130_fd_sc_hd__o41a_2 VGND X B1 A4 A3 A2 A1 VPWR VPB VNB
M$1 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=1610000U
M$3 VPWR B1 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=305000000000P AD=302500000000P PS=1610000U PD=1605000U
M$4 \$4 A4 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=302500000000P AD=177500000000P PS=1605000U PD=1355000U
M$5 \$14 A3 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=177500000000P AD=175000000000P PS=1355000U PD=1350000U
M$6 \$15 A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=175000000000P PS=1350000U PD=1350000U
M$7 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=410000000000P PS=1350000U PD=2820000U
M$8 \$4 B1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=208000000000P
+ AD=118625000000P PS=1940000U PD=1015000U
M$9 \$5 A4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=118625000000P AD=115375000000P PS=1015000U PD=1005000U
M$10 VGND A3 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=115375000000P AD=113750000000P PS=1005000U PD=1000000U
M$11 \$5 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=113750000000P PS=1000000U PD=1000000U
M$12 VGND A1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=113750000000P AD=266500000000P PS=1000000U PD=2120000U
M$13 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$14 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__o41a_2

.SUBCKT sky130_fd_sc_hd__decap_4 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1050000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1050000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__a31o_2 VPB X VPWR VGND A3 A2 A1 B1 VNB
M$1 VPWR \$10 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$10 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 VPWR A3 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 \$7 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=165000000000P PS=1270000U PD=1330000U
M$5 VPWR A1 \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=165000000000P PS=1330000U PD=1330000U
M$6 \$7 B1 \$10 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=320000000000P PS=1330000U PD=2640000U
M$7 VGND \$10 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=87750000000P PS=1820000U PD=920000U
M$8 X \$10 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$9 VGND A3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=87750000000P PS=920000U PD=920000U
M$10 \$13 A2 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=107250000000P PS=920000U PD=980000U
M$11 \$12 A1 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=126750000000P PS=980000U PD=1040000U
M$12 \$10 B1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=169000000000P PS=1040000U PD=1820000U
.ENDS sky130_fd_sc_hd__a31o_2

.SUBCKT sky130_fd_sc_hd__inv_2 VPB VGND VPWR Y A VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$3 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$4 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__mux2_1 VGND X A1 A0 S VPWR VPB VNB
M$1 VPWR S \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=158350000000P AD=76650000000P PS=1395000U PD=785000U
M$2 \$13 A0 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=76650000000P AD=193200000000P PS=785000U PD=1340000U
M$3 \$5 A1 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=193200000000P AD=44100000000P PS=1340000U PD=630000U
M$4 \$14 \$7 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=69300000000P PS=630000U PD=750000U
M$5 VPWR S \$7 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=69300000000P AD=117600000000P PS=750000U PD=1400000U
M$6 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=158350000000P PS=2520000U PD=1395000U
M$7 VGND S \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=112850000000P
+ AD=69300000000P PS=1045000U PD=750000U
M$8 \$8 A1 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=69300000000P
+ AD=99750000000P PS=750000U PD=895000U
M$9 \$5 A0 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=99750000000P
+ AD=69300000000P PS=895000U PD=750000U
M$10 \$9 \$7 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=69300000000P AD=144900000000P PS=750000U PD=1110000U
M$11 VGND S \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=144900000000P AD=109200000000P PS=1110000U PD=1360000U
M$12 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=112850000000P PS=1820000U PD=1045000U
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__o32a_2 VGND X A1 A2 A3 B2 B1 VPWR VPB VNB
M$1 VPWR \$5 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 X \$5 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=305000000000P PS=1270000U PD=1610000U
M$3 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=305000000000P AD=135000000000P PS=1610000U PD=1270000U
M$4 \$13 A2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=215000000000P PS=1270000U PD=1430000U
M$5 \$14 A3 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=215000000000P AD=135000000000P PS=1430000U PD=1270000U
M$6 \$5 B2 \$15 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=190000000000P PS=1270000U PD=1380000U
M$7 \$15 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=190000000000P AD=330000000000P PS=1380000U PD=2660000U
M$8 VGND \$5 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$5 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=198250000000P PS=920000U PD=1260000U
M$10 VGND A1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=198250000000P AD=87750000000P PS=1260000U PD=920000U
M$11 \$4 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=139750000000P PS=920000U PD=1080000U
M$12 VGND A3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=87750000000P PS=1080000U PD=920000U
M$13 \$4 B2 \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=123500000000P PS=920000U PD=1030000U
M$14 \$5 B1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=123500000000P AD=214500000000P PS=1030000U PD=1960000U
.ENDS sky130_fd_sc_hd__o32a_2

.SUBCKT sky130_fd_sc_hd__a32o_2 VGND X A1 A2 B2 B1 A3 VPWR VPB VNB
M$1 \$13 B2 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 \$4 B1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$13 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=215000000000P PS=1270000U PD=1430000U
M$4 VPWR A2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=215000000000P AD=135000000000P PS=1430000U PD=1270000U
M$5 \$13 A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$6 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$7 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=87750000000P PS=1820000U PD=920000U
M$9 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=209625000000P PS=920000U PD=1295000U
M$10 VGND B2 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=209625000000P AD=115375000000P PS=1295000U PD=1005000U
M$11 \$12 B1 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=115375000000P AD=107250000000P PS=1005000U PD=980000U
M$12 \$4 A1 \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=139750000000P PS=980000U PD=1080000U
M$13 \$11 A2 \$10 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=139750000000P AD=87750000000P PS=1080000U PD=920000U
M$14 \$10 A3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=87750000000P AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__a32o_2

.SUBCKT sky130_fd_sc_hd__clkbuf_1 VPB X VGND VPWR A VNB
M$1 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR A \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND A \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__o21ai_2 VPB A1 VGND A2 Y VPWR B1 VNB
M$1 VPWR A1 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 \$5 A2 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 Y A2 \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=175000000000P PS=1280000U PD=1350000U
M$4 \$5 A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=175000000000P AD=160000000000P PS=1350000U PD=1320000U
M$5 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=160000000000P AD=140000000000P PS=1320000U PD=1280000U
M$6 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$7 \$3 A1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=172250000000P AD=91000000000P PS=1830000U PD=930000U
M$8 VGND A2 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$9 \$3 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=126750000000P PS=930000U PD=1040000U
M$10 VGND A1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=126750000000P AD=91000000000P PS=1040000U PD=930000U
M$11 \$3 B1 Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=91000000000P PS=930000U PD=930000U
M$12 Y B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=91000000000P
+ AD=172250000000P PS=930000U PD=1830000U
.ENDS sky130_fd_sc_hd__o21ai_2

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__decap_6 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=1970000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=1970000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__nor2_2 VPB VGND A VPWR Y B VNB
M$1 \$4 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=280000000000P AD=135000000000P PS=2560000U PD=1270000U
M$2 VPWR A \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$3 \$4 B Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$4 Y B \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=182000000000P
+ AD=87750000000P PS=1860000U PD=920000U
M$6 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$7 VGND B Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=87750000000P PS=920000U PD=920000U
M$8 Y B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__nor2_2

.SUBCKT sky130_fd_sc_hd__decap_12 VPB VPWR VGND VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=4730000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=4730000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__fill_2 VPB VGND VPWR VNB
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__diode_2 VPB DIODE VPWR VGND VNB
D$1 DIODE VNB sky130_fd_pr__diode_pw2nd_05v5 A=434700000000P P=2640000U
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__clkinv_8 VGND Y A VPWR VPB VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=137500000000P PS=1270000U PD=1275000U
M$3 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=137500000000P AD=135000000000P PS=1275000U PD=1270000U
M$4 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$5 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$6 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$8 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$9 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$10 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$11 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$12 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$13 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=58800000000P PS=1370000U PD=700000U
M$14 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$15 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$16 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$17 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$18 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$19 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=58800000000P PS=700000U PD=700000U
M$20 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=111300000000P PS=700000U PD=1370000U
.ENDS sky130_fd_sc_hd__clkinv_8

.SUBCKT sky130_fd_sc_hd__clkinv_2 VPB Y A VPWR VGND VNB
M$1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=265000000000P AD=140000000000P PS=2530000U PD=1280000U
M$2 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=140000000000P PS=1280000U PD=1280000U
M$3 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=140000000000P AD=265000000000P PS=1280000U PD=2530000U
M$4 VGND A Y VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=111300000000P
+ AD=58800000000P PS=1370000U PD=700000U
M$5 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=58800000000P
+ AD=109200000000P PS=700000U PD=1360000U
.ENDS sky130_fd_sc_hd__clkinv_2

.SUBCKT sky130_fd_sc_hd__clkinv_1 VPB VPWR VGND Y A VNB
M$1 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=113400000000P PS=2200000U PD=1110000U
M$2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=113400000000P AD=235200000000P PS=1110000U PD=2240000U
M$3 Y A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=119700000000P PS=1360000U PD=1410000U
.ENDS sky130_fd_sc_hd__clkinv_1

.SUBCKT sky130_fd_sc_hd__decap_3 VPB VGND VPWR VNB
M$1 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=590000U W=870000U
+ AS=226200000000P AD=226200000000P PS=2260000U PD=2260000U
M$2 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 L=590000U W=550000U
+ AS=143000000000P AD=143000000000P PS=1620000U PD=1620000U
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__a221o_2 VGND B1 A1 X C1 B2 A2 VPWR VPB VNB
M$1 VPWR A1 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=165000000000P PS=2520000U PD=1330000U
M$2 \$13 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=157500000000P PS=1330000U PD=1315000U
M$3 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=135000000000P PS=1315000U PD=1270000U
M$4 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=285000000000P PS=1270000U PD=2570000U
M$5 \$3 C1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$12 B2 \$13 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=135000000000P PS=1270000U PD=1270000U
M$7 \$13 B1 \$12 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$8 \$3 A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=107250000000P PS=1820000U PD=980000U
M$9 \$8 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=102375000000P PS=980000U PD=965000U
M$10 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=102375000000P AD=87750000000P PS=965000U PD=920000U
M$11 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=185250000000P PS=920000U PD=1870000U
M$12 \$3 C1 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=107250000000P PS=1820000U PD=980000U
M$13 VGND B2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=68250000000P PS=980000U PD=860000U
M$14 \$7 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=68250000000P
+ AD=169000000000P PS=860000U PD=1820000U
.ENDS sky130_fd_sc_hd__a221o_2

.SUBCKT sky130_fd_sc_hd__or2_2 VPB X VPWR VGND B A VNB
M$1 \$4 B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=44100000000P PS=1360000U PD=630000U
M$2 \$9 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=44100000000P AD=155750000000P PS=630000U PD=1355000U
M$3 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=155750000000P AD=135000000000P PS=1355000U PD=1270000U
M$4 X \$4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$5 VGND B \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=109200000000P
+ AD=56700000000P PS=1360000U PD=690000U
M$6 \$4 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U AS=56700000000P
+ AD=106750000000P PS=690000U PD=1005000U
M$7 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=106750000000P
+ AD=87750000000P PS=1005000U PD=920000U
M$8 X \$4 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
.ENDS sky130_fd_sc_hd__or2_2

.SUBCKT sky130_fd_sc_hd__fill_1 VPB VGND VPWR VNB
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__a22o_2 VGND B1 A1 X B2 A2 VPWR VPB VNB
M$1 VPWR A1 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=165000000000P PS=2520000U PD=1330000U
M$2 \$11 A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=165000000000P AD=157500000000P PS=1330000U PD=1315000U
M$3 VPWR \$3 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=157500000000P AD=135000000000P PS=1315000U PD=1270000U
M$4 X \$3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=270000000000P PS=1270000U PD=2540000U
M$5 \$3 B2 \$11 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=260000000000P AD=135000000000P PS=2520000U PD=1270000U
M$6 \$11 B1 \$3 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$7 \$3 A1 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=169000000000P
+ AD=107250000000P PS=1820000U PD=980000U
M$8 \$8 A2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=107250000000P AD=102375000000P PS=980000U PD=965000U
M$9 VGND \$3 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=102375000000P
+ AD=87750000000P PS=965000U PD=920000U
M$10 X \$3 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=175500000000P PS=920000U PD=1840000U
M$11 VGND B2 \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=169000000000P AD=74750000000P PS=1820000U PD=880000U
M$12 \$7 B1 \$3 VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=74750000000P
+ AD=169000000000P PS=880000U PD=1820000U
.ENDS sky130_fd_sc_hd__a22o_2

.SUBCKT sky130_fd_sc_hd__o2bb2a_2 VGND X A2_N A1_N B2 B1 VPWR VPB VNB
M$1 VPWR \$8 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=285000000000P AD=135000000000P PS=2570000U PD=1270000U
M$2 X \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=154000000000P PS=1270000U PD=1335000U
M$3 VPWR A1_N \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=154000000000P AD=173000000000P PS=1335000U PD=1400000U
M$4 \$5 A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=173000000000P AD=227200000000P PS=1400000U PD=1350000U
M$5 VPWR \$5 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=227200000000P AD=92800000000P PS=1350000U PD=930000U
M$6 \$8 B2 \$14 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=92800000000P AD=86400000000P PS=930000U PD=910000U
M$7 \$14 B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$8 VGND A1_N \$7 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=98625000000P AD=66150000000P PS=980000U PD=735000U
M$9 \$7 A2_N \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66150000000P AD=109200000000P PS=735000U PD=1360000U
M$10 VGND \$8 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=185250000000P AD=87750000000P PS=1870000U PD=920000U
M$11 X \$8 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=98625000000P PS=920000U PD=980000U
M$12 \$8 \$5 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$13 \$6 B2 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=56700000000P PS=690000U PD=690000U
M$14 VGND B1 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
.ENDS sky130_fd_sc_hd__o2bb2a_2

.SUBCKT sky130_fd_sc_hd__buf_1 VPB X VGND VPWR A VNB
M$1 \$4 A VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=205400000000P AD=114550000000P PS=2100000U PD=1080000U
M$2 VPWR \$4 X VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=790000U
+ AS=114550000000P AD=205400000000P PS=1080000U PD=2100000U
M$3 \$4 A VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=135200000000P
+ AD=75400000000P PS=1560000U PD=810000U
M$4 VGND \$4 X VNB sky130_fd_pr__nfet_01v8 L=150000U W=520000U AS=75400000000P
+ AD=135200000000P PS=810000U PD=1560000U
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__dfrtp_2 VGND RESET_B Q CLK D VPWR VPB VNB
M$1 VPWR \$9 Q VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=301200000000P AD=135000000000P PS=2660000U PD=1270000U
M$2 Q \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=1000000U
+ AS=135000000000P AD=260000000000P PS=1270000U PD=2520000U
M$3 VPWR \$6 \$17 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=840000U
+ AS=218400000000P AD=129150000000P PS=2200000U PD=1185000U
M$4 \$17 \$3 \$8 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=129150000000P AD=58800000000P PS=1185000U PD=700000U
M$5 \$8 \$4 \$21 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=58800000000P AD=56700000000P PS=700000U PD=690000U
M$6 \$21 \$9 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=81900000000P PS=690000U PD=810000U
M$7 VPWR RESET_B \$9 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=81900000000P AD=56700000000P PS=810000U PD=690000U
M$8 \$9 \$8 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=56700000000P AD=113400000000P PS=690000U PD=1380000U
M$9 VPWR D \$5 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=109200000000P AD=65100000000P PS=1360000U PD=730000U
M$10 \$5 \$4 \$6 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=65100000000P AD=72450000000P PS=730000U PD=765000U
M$11 \$6 \$3 \$20 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=72450000000P AD=115500000000P PS=765000U PD=970000U
M$12 \$20 \$17 VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=115500000000P AD=70350000000P PS=970000U PD=755000U
M$13 VPWR RESET_B \$20 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=420000U
+ AS=70350000000P AD=109200000000P PS=755000U PD=1360000U
M$14 \$3 CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=166400000000P AD=86400000000P PS=1800000U PD=910000U
M$15 VPWR \$3 \$4 VPB sky130_fd_pr__pfet_01v8_hvt L=150000U W=640000U
+ AS=86400000000P AD=166400000000P PS=910000U PD=1800000U
M$16 VGND \$9 Q VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U
+ AS=208700000000P AD=87750000000P PS=2020000U PD=920000U
M$17 Q \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=650000U AS=87750000000P
+ AD=169000000000P PS=920000U PD=1820000U
M$18 \$3 CLK VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=109200000000P AD=56700000000P PS=1360000U PD=690000U
M$19 VGND \$3 \$4 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=56700000000P AD=109200000000P PS=690000U PD=1360000U
M$20 \$5 \$3 \$6 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=66000000000P AD=59400000000P PS=745000U PD=690000U
M$21 \$6 \$4 \$12 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=59400000000P AD=140100000000P PS=690000U PD=1100000U
M$22 \$17 \$4 \$8 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=99900000000P AD=71100000000P PS=985000U PD=755000U
M$23 \$8 \$3 \$13 VNB sky130_fd_pr__nfet_01v8 L=150000U W=360000U
+ AS=71100000000P AD=66900000000P PS=755000U PD=750000U
M$24 VGND D \$5 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=220500000000P AD=66000000000P PS=1890000U PD=745000U
M$25 \$12 \$17 \$14 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=140100000000P AD=44100000000P PS=1100000U PD=630000U
M$26 \$14 RESET_B VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=44100000000P AD=134600000000P PS=630000U PD=1150000U
M$27 \$13 \$9 VGND VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=66900000000P AD=124950000000P PS=750000U PD=1015000U
M$28 VGND RESET_B \$11 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=124950000000P AD=64050000000P PS=1015000U PD=725000U
M$29 \$11 \$8 \$9 VNB sky130_fd_pr__nfet_01v8 L=150000U W=420000U
+ AS=64050000000P AD=109200000000P PS=725000U PD=1360000U
M$30 VGND \$6 \$17 VNB sky130_fd_pr__nfet_01v8 L=150000U W=640000U
+ AS=134600000000P AD=99900000000P PS=1150000U PD=985000U
.ENDS sky130_fd_sc_hd__dfrtp_2
