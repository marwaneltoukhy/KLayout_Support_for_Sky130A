*SPICE netlist created from verilog structural netlist module mprj_logic_high by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /home/marwan/klayout_lvs/lvs/test_cases/mprj_logic_high/sky130_fd_sc_hd.spice

.subckt mprj_logic_high vccd1 vssd1 HI[0] HI[1] HI[2] HI[3] HI[4]
+ HI[5] HI[6] HI[7] HI[8] HI[9] HI[10] HI[11] HI[12]
+ HI[13] HI[14] HI[15] HI[16] HI[17] HI[18] HI[19] HI[20]
+ HI[21] HI[22] HI[23] HI[24] HI[25] HI[26] HI[27] HI[28]
+ HI[29] HI[30] HI[31] HI[32] HI[33] HI[34] HI[35] HI[36]
+ HI[37] HI[38] HI[39] HI[40] HI[41] HI[42] HI[43] HI[44]
+ HI[45] HI[46] HI[47] HI[48] HI[49] HI[50] HI[51] HI[52]
+ HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59] HI[60]
+ HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68]
+ HI[69] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76]
+ HI[77] HI[78] HI[79] HI[80] HI[81] HI[82] HI[83] HI[84]
+ HI[85] HI[86] HI[87] HI[88] HI[89] HI[90] HI[91] HI[92]
+ HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[100]
+ HI[101] HI[102] HI[103] HI[104] HI[105] HI[106] HI[107] HI[108]
+ HI[109] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[120] HI[121] HI[122] HI[123] HI[124]
+ HI[125] HI[126] HI[127] HI[128] HI[129] HI[130] HI[131] HI[132]
+ HI[133] HI[134] HI[135] HI[136] HI[137] HI[138] HI[139] HI[140]
+ HI[141] HI[142] HI[143] HI[144] HI[145] HI[146] HI[147] HI[148]
+ HI[149] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[160] HI[161] HI[162] HI[163] HI[164]
+ HI[165] HI[166] HI[167] HI[168] HI[169] HI[170] HI[171] HI[172]
+ HI[173] HI[174] HI[175] HI[176] HI[177] HI[178] HI[179] HI[180]
+ HI[181] HI[182] HI[183] HI[184] HI[185] HI[186] HI[187] HI[188]
+ HI[189] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[200] HI[201] HI[202] HI[203] HI[204]
+ HI[205] HI[206] HI[207] HI[208] HI[209] HI[210] HI[211] HI[212]
+ HI[213] HI[214] HI[215] HI[216] HI[217] HI[218] HI[219] HI[220]
+ HI[221] HI[222] HI[223] HI[224] HI[225] HI[226] HI[227] HI[228]
+ HI[229] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235] HI[236]
+ HI[237] HI[238] HI[239] HI[240] HI[241] HI[242] HI[243] HI[244]
+ HI[245] HI[246] HI[247] HI[248] HI[249] HI[250] HI[251] HI[252]
+ HI[253] HI[254] HI[255] HI[256] HI[257] HI[258] HI[259] HI[260]
+ HI[261] HI[262] HI[263] HI[264] HI[265] HI[266] HI[267] HI[268]
+ HI[269] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275] HI[276]
+ HI[277] HI[278] HI[279] HI[280] HI[281] HI[282] HI[283] HI[284]
+ HI[285] HI[286] HI[287] HI[288] HI[289] HI[290] HI[291] HI[292]
+ HI[293] HI[294] HI[295] HI[296] HI[297] HI[298] HI[299] HI[300]
+ HI[301] HI[302] HI[303] HI[304] HI[305] HI[306] HI[307] HI[308]
+ HI[309] HI[310] HI[311] HI[312] HI[313] HI[314] HI[315] HI[316]
+ HI[317] HI[318] HI[319] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[330] HI[331] HI[332]
+ HI[333] HI[334] HI[335] HI[336] HI[337] HI[338] HI[339] HI[340]
+ HI[341] HI[342] HI[343] HI[344] HI[345] HI[346] HI[347] HI[348]
+ HI[349] HI[350] HI[351] HI[352] HI[353] HI[354] HI[355] HI[356]
+ HI[357] HI[358] HI[359] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[370] HI[371] HI[372]
+ HI[373] HI[374] HI[375] HI[376] HI[377] HI[378] HI[379] HI[380]
+ HI[381] HI[382] HI[383] HI[384] HI[385] HI[386] HI[387] HI[388]
+ HI[389] HI[390] HI[391] HI[392] HI[393] HI[394] HI[395] HI[396]
+ HI[397] HI[398] HI[399] HI[400] HI[401] HI[402] HI[403] HI[404]
+ HI[405] HI[406] HI[407] HI[408] HI[409] HI[410] HI[411] HI[412]
+ HI[413] HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[420]
+ HI[421] HI[422] HI[423] HI[424] HI[425] HI[426] HI[427] HI[428]
+ HI[429] HI[430] HI[431] HI[432] HI[433] HI[434] HI[435] HI[436]
+ HI[437] HI[438] HI[439] HI[440] HI[441] HI[442] HI[443] HI[444]
+ HI[445] HI[446] HI[447] HI[448] HI[449] HI[450] HI[451] HI[452]
+ HI[453] HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[460]
+ HI[461] HI[462] 

XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_10 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_11 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_12 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_13 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_14 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_15 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_16 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_17 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_18 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_19 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_20 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_21 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_22 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_23 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_24 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_25 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_26 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_27 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_28 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_29 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_30 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_31 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_32 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_33 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_37 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_38 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_39 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_8 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_9 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X\insts[0]  vssd1 vssd1 vccd1 vccd1 HI[0] NC sky130_fd_sc_hd__conb_1
X\insts[100]  vssd1 vssd1 vccd1 vccd1 HI[100] NC sky130_fd_sc_hd__conb_1
X\insts[101]  vssd1 vssd1 vccd1 vccd1 HI[101] NC sky130_fd_sc_hd__conb_1
X\insts[102]  vssd1 vssd1 vccd1 vccd1 HI[102] NC sky130_fd_sc_hd__conb_1
X\insts[103]  vssd1 vssd1 vccd1 vccd1 HI[103] NC sky130_fd_sc_hd__conb_1
X\insts[104]  vssd1 vssd1 vccd1 vccd1 HI[104] NC sky130_fd_sc_hd__conb_1
X\insts[105]  vssd1 vssd1 vccd1 vccd1 HI[105] NC sky130_fd_sc_hd__conb_1
X\insts[106]  vssd1 vssd1 vccd1 vccd1 HI[106] NC sky130_fd_sc_hd__conb_1
X\insts[107]  vssd1 vssd1 vccd1 vccd1 HI[107] NC sky130_fd_sc_hd__conb_1
X\insts[108]  vssd1 vssd1 vccd1 vccd1 HI[108] NC sky130_fd_sc_hd__conb_1
X\insts[109]  vssd1 vssd1 vccd1 vccd1 HI[109] NC sky130_fd_sc_hd__conb_1
X\insts[10]  vssd1 vssd1 vccd1 vccd1 HI[10] NC sky130_fd_sc_hd__conb_1
X\insts[110]  vssd1 vssd1 vccd1 vccd1 HI[110] NC sky130_fd_sc_hd__conb_1
X\insts[111]  vssd1 vssd1 vccd1 vccd1 HI[111] NC sky130_fd_sc_hd__conb_1
X\insts[112]  vssd1 vssd1 vccd1 vccd1 HI[112] NC sky130_fd_sc_hd__conb_1
X\insts[113]  vssd1 vssd1 vccd1 vccd1 HI[113] NC sky130_fd_sc_hd__conb_1
X\insts[114]  vssd1 vssd1 vccd1 vccd1 HI[114] NC sky130_fd_sc_hd__conb_1
X\insts[115]  vssd1 vssd1 vccd1 vccd1 HI[115] NC sky130_fd_sc_hd__conb_1
X\insts[116]  vssd1 vssd1 vccd1 vccd1 HI[116] NC sky130_fd_sc_hd__conb_1
X\insts[117]  vssd1 vssd1 vccd1 vccd1 HI[117] NC sky130_fd_sc_hd__conb_1
X\insts[118]  vssd1 vssd1 vccd1 vccd1 HI[118] NC sky130_fd_sc_hd__conb_1
X\insts[119]  vssd1 vssd1 vccd1 vccd1 HI[119] NC sky130_fd_sc_hd__conb_1
X\insts[11]  vssd1 vssd1 vccd1 vccd1 HI[11] NC sky130_fd_sc_hd__conb_1
X\insts[120]  vssd1 vssd1 vccd1 vccd1 HI[120] NC sky130_fd_sc_hd__conb_1
X\insts[121]  vssd1 vssd1 vccd1 vccd1 HI[121] NC sky130_fd_sc_hd__conb_1
X\insts[122]  vssd1 vssd1 vccd1 vccd1 HI[122] NC sky130_fd_sc_hd__conb_1
X\insts[123]  vssd1 vssd1 vccd1 vccd1 HI[123] NC sky130_fd_sc_hd__conb_1
X\insts[124]  vssd1 vssd1 vccd1 vccd1 HI[124] NC sky130_fd_sc_hd__conb_1
X\insts[125]  vssd1 vssd1 vccd1 vccd1 HI[125] NC sky130_fd_sc_hd__conb_1
X\insts[126]  vssd1 vssd1 vccd1 vccd1 HI[126] NC sky130_fd_sc_hd__conb_1
X\insts[127]  vssd1 vssd1 vccd1 vccd1 HI[127] NC sky130_fd_sc_hd__conb_1
X\insts[128]  vssd1 vssd1 vccd1 vccd1 HI[128] NC sky130_fd_sc_hd__conb_1
X\insts[129]  vssd1 vssd1 vccd1 vccd1 HI[129] NC sky130_fd_sc_hd__conb_1
X\insts[12]  vssd1 vssd1 vccd1 vccd1 HI[12] NC sky130_fd_sc_hd__conb_1
X\insts[130]  vssd1 vssd1 vccd1 vccd1 HI[130] NC sky130_fd_sc_hd__conb_1
X\insts[131]  vssd1 vssd1 vccd1 vccd1 HI[131] NC sky130_fd_sc_hd__conb_1
X\insts[132]  vssd1 vssd1 vccd1 vccd1 HI[132] NC sky130_fd_sc_hd__conb_1
X\insts[133]  vssd1 vssd1 vccd1 vccd1 HI[133] NC sky130_fd_sc_hd__conb_1
X\insts[134]  vssd1 vssd1 vccd1 vccd1 HI[134] NC sky130_fd_sc_hd__conb_1
X\insts[135]  vssd1 vssd1 vccd1 vccd1 HI[135] NC sky130_fd_sc_hd__conb_1
X\insts[136]  vssd1 vssd1 vccd1 vccd1 HI[136] NC sky130_fd_sc_hd__conb_1
X\insts[137]  vssd1 vssd1 vccd1 vccd1 HI[137] NC sky130_fd_sc_hd__conb_1
X\insts[138]  vssd1 vssd1 vccd1 vccd1 HI[138] NC sky130_fd_sc_hd__conb_1
X\insts[139]  vssd1 vssd1 vccd1 vccd1 HI[139] NC sky130_fd_sc_hd__conb_1
X\insts[13]  vssd1 vssd1 vccd1 vccd1 HI[13] NC sky130_fd_sc_hd__conb_1
X\insts[140]  vssd1 vssd1 vccd1 vccd1 HI[140] NC sky130_fd_sc_hd__conb_1
X\insts[141]  vssd1 vssd1 vccd1 vccd1 HI[141] NC sky130_fd_sc_hd__conb_1
X\insts[142]  vssd1 vssd1 vccd1 vccd1 HI[142] NC sky130_fd_sc_hd__conb_1
X\insts[143]  vssd1 vssd1 vccd1 vccd1 HI[143] NC sky130_fd_sc_hd__conb_1
X\insts[144]  vssd1 vssd1 vccd1 vccd1 HI[144] NC sky130_fd_sc_hd__conb_1
X\insts[145]  vssd1 vssd1 vccd1 vccd1 HI[145] NC sky130_fd_sc_hd__conb_1
X\insts[146]  vssd1 vssd1 vccd1 vccd1 HI[146] NC sky130_fd_sc_hd__conb_1
X\insts[147]  vssd1 vssd1 vccd1 vccd1 HI[147] NC sky130_fd_sc_hd__conb_1
X\insts[148]  vssd1 vssd1 vccd1 vccd1 HI[148] NC sky130_fd_sc_hd__conb_1
X\insts[149]  vssd1 vssd1 vccd1 vccd1 HI[149] NC sky130_fd_sc_hd__conb_1
X\insts[14]  vssd1 vssd1 vccd1 vccd1 HI[14] NC sky130_fd_sc_hd__conb_1
X\insts[150]  vssd1 vssd1 vccd1 vccd1 HI[150] NC sky130_fd_sc_hd__conb_1
X\insts[151]  vssd1 vssd1 vccd1 vccd1 HI[151] NC sky130_fd_sc_hd__conb_1
X\insts[152]  vssd1 vssd1 vccd1 vccd1 HI[152] NC sky130_fd_sc_hd__conb_1
X\insts[153]  vssd1 vssd1 vccd1 vccd1 HI[153] NC sky130_fd_sc_hd__conb_1
X\insts[154]  vssd1 vssd1 vccd1 vccd1 HI[154] NC sky130_fd_sc_hd__conb_1
X\insts[155]  vssd1 vssd1 vccd1 vccd1 HI[155] NC sky130_fd_sc_hd__conb_1
X\insts[156]  vssd1 vssd1 vccd1 vccd1 HI[156] NC sky130_fd_sc_hd__conb_1
X\insts[157]  vssd1 vssd1 vccd1 vccd1 HI[157] NC sky130_fd_sc_hd__conb_1
X\insts[158]  vssd1 vssd1 vccd1 vccd1 HI[158] NC sky130_fd_sc_hd__conb_1
X\insts[159]  vssd1 vssd1 vccd1 vccd1 HI[159] NC sky130_fd_sc_hd__conb_1
X\insts[15]  vssd1 vssd1 vccd1 vccd1 HI[15] NC sky130_fd_sc_hd__conb_1
X\insts[160]  vssd1 vssd1 vccd1 vccd1 HI[160] NC sky130_fd_sc_hd__conb_1
X\insts[161]  vssd1 vssd1 vccd1 vccd1 HI[161] NC sky130_fd_sc_hd__conb_1
X\insts[162]  vssd1 vssd1 vccd1 vccd1 HI[162] NC sky130_fd_sc_hd__conb_1
X\insts[163]  vssd1 vssd1 vccd1 vccd1 HI[163] NC sky130_fd_sc_hd__conb_1
X\insts[164]  vssd1 vssd1 vccd1 vccd1 HI[164] NC sky130_fd_sc_hd__conb_1
X\insts[165]  vssd1 vssd1 vccd1 vccd1 HI[165] NC sky130_fd_sc_hd__conb_1
X\insts[166]  vssd1 vssd1 vccd1 vccd1 HI[166] NC sky130_fd_sc_hd__conb_1
X\insts[167]  vssd1 vssd1 vccd1 vccd1 HI[167] NC sky130_fd_sc_hd__conb_1
X\insts[168]  vssd1 vssd1 vccd1 vccd1 HI[168] NC sky130_fd_sc_hd__conb_1
X\insts[169]  vssd1 vssd1 vccd1 vccd1 HI[169] NC sky130_fd_sc_hd__conb_1
X\insts[16]  vssd1 vssd1 vccd1 vccd1 HI[16] NC sky130_fd_sc_hd__conb_1
X\insts[170]  vssd1 vssd1 vccd1 vccd1 HI[170] NC sky130_fd_sc_hd__conb_1
X\insts[171]  vssd1 vssd1 vccd1 vccd1 HI[171] NC sky130_fd_sc_hd__conb_1
X\insts[172]  vssd1 vssd1 vccd1 vccd1 HI[172] NC sky130_fd_sc_hd__conb_1
X\insts[173]  vssd1 vssd1 vccd1 vccd1 HI[173] NC sky130_fd_sc_hd__conb_1
X\insts[174]  vssd1 vssd1 vccd1 vccd1 HI[174] NC sky130_fd_sc_hd__conb_1
X\insts[175]  vssd1 vssd1 vccd1 vccd1 HI[175] NC sky130_fd_sc_hd__conb_1
X\insts[176]  vssd1 vssd1 vccd1 vccd1 HI[176] NC sky130_fd_sc_hd__conb_1
X\insts[177]  vssd1 vssd1 vccd1 vccd1 HI[177] NC sky130_fd_sc_hd__conb_1
X\insts[178]  vssd1 vssd1 vccd1 vccd1 HI[178] NC sky130_fd_sc_hd__conb_1
X\insts[179]  vssd1 vssd1 vccd1 vccd1 HI[179] NC sky130_fd_sc_hd__conb_1
X\insts[17]  vssd1 vssd1 vccd1 vccd1 HI[17] NC sky130_fd_sc_hd__conb_1
X\insts[180]  vssd1 vssd1 vccd1 vccd1 HI[180] NC sky130_fd_sc_hd__conb_1
X\insts[181]  vssd1 vssd1 vccd1 vccd1 HI[181] NC sky130_fd_sc_hd__conb_1
X\insts[182]  vssd1 vssd1 vccd1 vccd1 HI[182] NC sky130_fd_sc_hd__conb_1
X\insts[183]  vssd1 vssd1 vccd1 vccd1 HI[183] NC sky130_fd_sc_hd__conb_1
X\insts[184]  vssd1 vssd1 vccd1 vccd1 HI[184] NC sky130_fd_sc_hd__conb_1
X\insts[185]  vssd1 vssd1 vccd1 vccd1 HI[185] NC sky130_fd_sc_hd__conb_1
X\insts[186]  vssd1 vssd1 vccd1 vccd1 HI[186] NC sky130_fd_sc_hd__conb_1
X\insts[187]  vssd1 vssd1 vccd1 vccd1 HI[187] NC sky130_fd_sc_hd__conb_1
X\insts[188]  vssd1 vssd1 vccd1 vccd1 HI[188] NC sky130_fd_sc_hd__conb_1
X\insts[189]  vssd1 vssd1 vccd1 vccd1 HI[189] NC sky130_fd_sc_hd__conb_1
X\insts[18]  vssd1 vssd1 vccd1 vccd1 HI[18] NC sky130_fd_sc_hd__conb_1
X\insts[190]  vssd1 vssd1 vccd1 vccd1 HI[190] NC sky130_fd_sc_hd__conb_1
X\insts[191]  vssd1 vssd1 vccd1 vccd1 HI[191] NC sky130_fd_sc_hd__conb_1
X\insts[192]  vssd1 vssd1 vccd1 vccd1 HI[192] NC sky130_fd_sc_hd__conb_1
X\insts[193]  vssd1 vssd1 vccd1 vccd1 HI[193] NC sky130_fd_sc_hd__conb_1
X\insts[194]  vssd1 vssd1 vccd1 vccd1 HI[194] NC sky130_fd_sc_hd__conb_1
X\insts[195]  vssd1 vssd1 vccd1 vccd1 HI[195] NC sky130_fd_sc_hd__conb_1
X\insts[196]  vssd1 vssd1 vccd1 vccd1 HI[196] NC sky130_fd_sc_hd__conb_1
X\insts[197]  vssd1 vssd1 vccd1 vccd1 HI[197] NC sky130_fd_sc_hd__conb_1
X\insts[198]  vssd1 vssd1 vccd1 vccd1 HI[198] NC sky130_fd_sc_hd__conb_1
X\insts[199]  vssd1 vssd1 vccd1 vccd1 HI[199] NC sky130_fd_sc_hd__conb_1
X\insts[19]  vssd1 vssd1 vccd1 vccd1 HI[19] NC sky130_fd_sc_hd__conb_1
X\insts[1]  vssd1 vssd1 vccd1 vccd1 HI[1] NC sky130_fd_sc_hd__conb_1
X\insts[200]  vssd1 vssd1 vccd1 vccd1 HI[200] NC sky130_fd_sc_hd__conb_1
X\insts[201]  vssd1 vssd1 vccd1 vccd1 HI[201] NC sky130_fd_sc_hd__conb_1
X\insts[202]  vssd1 vssd1 vccd1 vccd1 HI[202] NC sky130_fd_sc_hd__conb_1
X\insts[203]  vssd1 vssd1 vccd1 vccd1 HI[203] NC sky130_fd_sc_hd__conb_1
X\insts[204]  vssd1 vssd1 vccd1 vccd1 HI[204] NC sky130_fd_sc_hd__conb_1
X\insts[205]  vssd1 vssd1 vccd1 vccd1 HI[205] NC sky130_fd_sc_hd__conb_1
X\insts[206]  vssd1 vssd1 vccd1 vccd1 HI[206] NC sky130_fd_sc_hd__conb_1
X\insts[207]  vssd1 vssd1 vccd1 vccd1 HI[207] NC sky130_fd_sc_hd__conb_1
X\insts[208]  vssd1 vssd1 vccd1 vccd1 HI[208] NC sky130_fd_sc_hd__conb_1
X\insts[209]  vssd1 vssd1 vccd1 vccd1 HI[209] NC sky130_fd_sc_hd__conb_1
X\insts[20]  vssd1 vssd1 vccd1 vccd1 HI[20] NC sky130_fd_sc_hd__conb_1
X\insts[210]  vssd1 vssd1 vccd1 vccd1 HI[210] NC sky130_fd_sc_hd__conb_1
X\insts[211]  vssd1 vssd1 vccd1 vccd1 HI[211] NC sky130_fd_sc_hd__conb_1
X\insts[212]  vssd1 vssd1 vccd1 vccd1 HI[212] NC sky130_fd_sc_hd__conb_1
X\insts[213]  vssd1 vssd1 vccd1 vccd1 HI[213] NC sky130_fd_sc_hd__conb_1
X\insts[214]  vssd1 vssd1 vccd1 vccd1 HI[214] NC sky130_fd_sc_hd__conb_1
X\insts[215]  vssd1 vssd1 vccd1 vccd1 HI[215] NC sky130_fd_sc_hd__conb_1
X\insts[216]  vssd1 vssd1 vccd1 vccd1 HI[216] NC sky130_fd_sc_hd__conb_1
X\insts[217]  vssd1 vssd1 vccd1 vccd1 HI[217] NC sky130_fd_sc_hd__conb_1
X\insts[218]  vssd1 vssd1 vccd1 vccd1 HI[218] NC sky130_fd_sc_hd__conb_1
X\insts[219]  vssd1 vssd1 vccd1 vccd1 HI[219] NC sky130_fd_sc_hd__conb_1
X\insts[21]  vssd1 vssd1 vccd1 vccd1 HI[21] NC sky130_fd_sc_hd__conb_1
X\insts[220]  vssd1 vssd1 vccd1 vccd1 HI[220] NC sky130_fd_sc_hd__conb_1
X\insts[221]  vssd1 vssd1 vccd1 vccd1 HI[221] NC sky130_fd_sc_hd__conb_1
X\insts[222]  vssd1 vssd1 vccd1 vccd1 HI[222] NC sky130_fd_sc_hd__conb_1
X\insts[223]  vssd1 vssd1 vccd1 vccd1 HI[223] NC sky130_fd_sc_hd__conb_1
X\insts[224]  vssd1 vssd1 vccd1 vccd1 HI[224] NC sky130_fd_sc_hd__conb_1
X\insts[225]  vssd1 vssd1 vccd1 vccd1 HI[225] NC sky130_fd_sc_hd__conb_1
X\insts[226]  vssd1 vssd1 vccd1 vccd1 HI[226] NC sky130_fd_sc_hd__conb_1
X\insts[227]  vssd1 vssd1 vccd1 vccd1 HI[227] NC sky130_fd_sc_hd__conb_1
X\insts[228]  vssd1 vssd1 vccd1 vccd1 HI[228] NC sky130_fd_sc_hd__conb_1
X\insts[229]  vssd1 vssd1 vccd1 vccd1 HI[229] NC sky130_fd_sc_hd__conb_1
X\insts[22]  vssd1 vssd1 vccd1 vccd1 HI[22] NC sky130_fd_sc_hd__conb_1
X\insts[230]  vssd1 vssd1 vccd1 vccd1 HI[230] NC sky130_fd_sc_hd__conb_1
X\insts[231]  vssd1 vssd1 vccd1 vccd1 HI[231] NC sky130_fd_sc_hd__conb_1
X\insts[232]  vssd1 vssd1 vccd1 vccd1 HI[232] NC sky130_fd_sc_hd__conb_1
X\insts[233]  vssd1 vssd1 vccd1 vccd1 HI[233] NC sky130_fd_sc_hd__conb_1
X\insts[234]  vssd1 vssd1 vccd1 vccd1 HI[234] NC sky130_fd_sc_hd__conb_1
X\insts[235]  vssd1 vssd1 vccd1 vccd1 HI[235] NC sky130_fd_sc_hd__conb_1
X\insts[236]  vssd1 vssd1 vccd1 vccd1 HI[236] NC sky130_fd_sc_hd__conb_1
X\insts[237]  vssd1 vssd1 vccd1 vccd1 HI[237] NC sky130_fd_sc_hd__conb_1
X\insts[238]  vssd1 vssd1 vccd1 vccd1 HI[238] NC sky130_fd_sc_hd__conb_1
X\insts[239]  vssd1 vssd1 vccd1 vccd1 HI[239] NC sky130_fd_sc_hd__conb_1
X\insts[23]  vssd1 vssd1 vccd1 vccd1 HI[23] NC sky130_fd_sc_hd__conb_1
X\insts[240]  vssd1 vssd1 vccd1 vccd1 HI[240] NC sky130_fd_sc_hd__conb_1
X\insts[241]  vssd1 vssd1 vccd1 vccd1 HI[241] NC sky130_fd_sc_hd__conb_1
X\insts[242]  vssd1 vssd1 vccd1 vccd1 HI[242] NC sky130_fd_sc_hd__conb_1
X\insts[243]  vssd1 vssd1 vccd1 vccd1 HI[243] NC sky130_fd_sc_hd__conb_1
X\insts[244]  vssd1 vssd1 vccd1 vccd1 HI[244] NC sky130_fd_sc_hd__conb_1
X\insts[245]  vssd1 vssd1 vccd1 vccd1 HI[245] NC sky130_fd_sc_hd__conb_1
X\insts[246]  vssd1 vssd1 vccd1 vccd1 HI[246] NC sky130_fd_sc_hd__conb_1
X\insts[247]  vssd1 vssd1 vccd1 vccd1 HI[247] NC sky130_fd_sc_hd__conb_1
X\insts[248]  vssd1 vssd1 vccd1 vccd1 HI[248] NC sky130_fd_sc_hd__conb_1
X\insts[249]  vssd1 vssd1 vccd1 vccd1 HI[249] NC sky130_fd_sc_hd__conb_1
X\insts[24]  vssd1 vssd1 vccd1 vccd1 HI[24] NC sky130_fd_sc_hd__conb_1
X\insts[250]  vssd1 vssd1 vccd1 vccd1 HI[250] NC sky130_fd_sc_hd__conb_1
X\insts[251]  vssd1 vssd1 vccd1 vccd1 HI[251] NC sky130_fd_sc_hd__conb_1
X\insts[252]  vssd1 vssd1 vccd1 vccd1 HI[252] NC sky130_fd_sc_hd__conb_1
X\insts[253]  vssd1 vssd1 vccd1 vccd1 HI[253] NC sky130_fd_sc_hd__conb_1
X\insts[254]  vssd1 vssd1 vccd1 vccd1 HI[254] NC sky130_fd_sc_hd__conb_1
X\insts[255]  vssd1 vssd1 vccd1 vccd1 HI[255] NC sky130_fd_sc_hd__conb_1
X\insts[256]  vssd1 vssd1 vccd1 vccd1 HI[256] NC sky130_fd_sc_hd__conb_1
X\insts[257]  vssd1 vssd1 vccd1 vccd1 HI[257] NC sky130_fd_sc_hd__conb_1
X\insts[258]  vssd1 vssd1 vccd1 vccd1 HI[258] NC sky130_fd_sc_hd__conb_1
X\insts[259]  vssd1 vssd1 vccd1 vccd1 HI[259] NC sky130_fd_sc_hd__conb_1
X\insts[25]  vssd1 vssd1 vccd1 vccd1 HI[25] NC sky130_fd_sc_hd__conb_1
X\insts[260]  vssd1 vssd1 vccd1 vccd1 HI[260] NC sky130_fd_sc_hd__conb_1
X\insts[261]  vssd1 vssd1 vccd1 vccd1 HI[261] NC sky130_fd_sc_hd__conb_1
X\insts[262]  vssd1 vssd1 vccd1 vccd1 HI[262] NC sky130_fd_sc_hd__conb_1
X\insts[263]  vssd1 vssd1 vccd1 vccd1 HI[263] NC sky130_fd_sc_hd__conb_1
X\insts[264]  vssd1 vssd1 vccd1 vccd1 HI[264] NC sky130_fd_sc_hd__conb_1
X\insts[265]  vssd1 vssd1 vccd1 vccd1 HI[265] NC sky130_fd_sc_hd__conb_1
X\insts[266]  vssd1 vssd1 vccd1 vccd1 HI[266] NC sky130_fd_sc_hd__conb_1
X\insts[267]  vssd1 vssd1 vccd1 vccd1 HI[267] NC sky130_fd_sc_hd__conb_1
X\insts[268]  vssd1 vssd1 vccd1 vccd1 HI[268] NC sky130_fd_sc_hd__conb_1
X\insts[269]  vssd1 vssd1 vccd1 vccd1 HI[269] NC sky130_fd_sc_hd__conb_1
X\insts[26]  vssd1 vssd1 vccd1 vccd1 HI[26] NC sky130_fd_sc_hd__conb_1
X\insts[270]  vssd1 vssd1 vccd1 vccd1 HI[270] NC sky130_fd_sc_hd__conb_1
X\insts[271]  vssd1 vssd1 vccd1 vccd1 HI[271] NC sky130_fd_sc_hd__conb_1
X\insts[272]  vssd1 vssd1 vccd1 vccd1 HI[272] NC sky130_fd_sc_hd__conb_1
X\insts[273]  vssd1 vssd1 vccd1 vccd1 HI[273] NC sky130_fd_sc_hd__conb_1
X\insts[274]  vssd1 vssd1 vccd1 vccd1 HI[274] NC sky130_fd_sc_hd__conb_1
X\insts[275]  vssd1 vssd1 vccd1 vccd1 HI[275] NC sky130_fd_sc_hd__conb_1
X\insts[276]  vssd1 vssd1 vccd1 vccd1 HI[276] NC sky130_fd_sc_hd__conb_1
X\insts[277]  vssd1 vssd1 vccd1 vccd1 HI[277] NC sky130_fd_sc_hd__conb_1
X\insts[278]  vssd1 vssd1 vccd1 vccd1 HI[278] NC sky130_fd_sc_hd__conb_1
X\insts[279]  vssd1 vssd1 vccd1 vccd1 HI[279] NC sky130_fd_sc_hd__conb_1
X\insts[27]  vssd1 vssd1 vccd1 vccd1 HI[27] NC sky130_fd_sc_hd__conb_1
X\insts[280]  vssd1 vssd1 vccd1 vccd1 HI[280] NC sky130_fd_sc_hd__conb_1
X\insts[281]  vssd1 vssd1 vccd1 vccd1 HI[281] NC sky130_fd_sc_hd__conb_1
X\insts[282]  vssd1 vssd1 vccd1 vccd1 HI[282] NC sky130_fd_sc_hd__conb_1
X\insts[283]  vssd1 vssd1 vccd1 vccd1 HI[283] NC sky130_fd_sc_hd__conb_1
X\insts[284]  vssd1 vssd1 vccd1 vccd1 HI[284] NC sky130_fd_sc_hd__conb_1
X\insts[285]  vssd1 vssd1 vccd1 vccd1 HI[285] NC sky130_fd_sc_hd__conb_1
X\insts[286]  vssd1 vssd1 vccd1 vccd1 HI[286] NC sky130_fd_sc_hd__conb_1
X\insts[287]  vssd1 vssd1 vccd1 vccd1 HI[287] NC sky130_fd_sc_hd__conb_1
X\insts[288]  vssd1 vssd1 vccd1 vccd1 HI[288] NC sky130_fd_sc_hd__conb_1
X\insts[289]  vssd1 vssd1 vccd1 vccd1 HI[289] NC sky130_fd_sc_hd__conb_1
X\insts[28]  vssd1 vssd1 vccd1 vccd1 HI[28] NC sky130_fd_sc_hd__conb_1
X\insts[290]  vssd1 vssd1 vccd1 vccd1 HI[290] NC sky130_fd_sc_hd__conb_1
X\insts[291]  vssd1 vssd1 vccd1 vccd1 HI[291] NC sky130_fd_sc_hd__conb_1
X\insts[292]  vssd1 vssd1 vccd1 vccd1 HI[292] NC sky130_fd_sc_hd__conb_1
X\insts[293]  vssd1 vssd1 vccd1 vccd1 HI[293] NC sky130_fd_sc_hd__conb_1
X\insts[294]  vssd1 vssd1 vccd1 vccd1 HI[294] NC sky130_fd_sc_hd__conb_1
X\insts[295]  vssd1 vssd1 vccd1 vccd1 HI[295] NC sky130_fd_sc_hd__conb_1
X\insts[296]  vssd1 vssd1 vccd1 vccd1 HI[296] NC sky130_fd_sc_hd__conb_1
X\insts[297]  vssd1 vssd1 vccd1 vccd1 HI[297] NC sky130_fd_sc_hd__conb_1
X\insts[298]  vssd1 vssd1 vccd1 vccd1 HI[298] NC sky130_fd_sc_hd__conb_1
X\insts[299]  vssd1 vssd1 vccd1 vccd1 HI[299] NC sky130_fd_sc_hd__conb_1
X\insts[29]  vssd1 vssd1 vccd1 vccd1 HI[29] NC sky130_fd_sc_hd__conb_1
X\insts[2]  vssd1 vssd1 vccd1 vccd1 HI[2] NC sky130_fd_sc_hd__conb_1
X\insts[300]  vssd1 vssd1 vccd1 vccd1 HI[300] NC sky130_fd_sc_hd__conb_1
X\insts[301]  vssd1 vssd1 vccd1 vccd1 HI[301] NC sky130_fd_sc_hd__conb_1
X\insts[302]  vssd1 vssd1 vccd1 vccd1 HI[302] NC sky130_fd_sc_hd__conb_1
X\insts[303]  vssd1 vssd1 vccd1 vccd1 HI[303] NC sky130_fd_sc_hd__conb_1
X\insts[304]  vssd1 vssd1 vccd1 vccd1 HI[304] NC sky130_fd_sc_hd__conb_1
X\insts[305]  vssd1 vssd1 vccd1 vccd1 HI[305] NC sky130_fd_sc_hd__conb_1
X\insts[306]  vssd1 vssd1 vccd1 vccd1 HI[306] NC sky130_fd_sc_hd__conb_1
X\insts[307]  vssd1 vssd1 vccd1 vccd1 HI[307] NC sky130_fd_sc_hd__conb_1
X\insts[308]  vssd1 vssd1 vccd1 vccd1 HI[308] NC sky130_fd_sc_hd__conb_1
X\insts[309]  vssd1 vssd1 vccd1 vccd1 HI[309] NC sky130_fd_sc_hd__conb_1
X\insts[30]  vssd1 vssd1 vccd1 vccd1 HI[30] NC sky130_fd_sc_hd__conb_1
X\insts[310]  vssd1 vssd1 vccd1 vccd1 HI[310] NC sky130_fd_sc_hd__conb_1
X\insts[311]  vssd1 vssd1 vccd1 vccd1 HI[311] NC sky130_fd_sc_hd__conb_1
X\insts[312]  vssd1 vssd1 vccd1 vccd1 HI[312] NC sky130_fd_sc_hd__conb_1
X\insts[313]  vssd1 vssd1 vccd1 vccd1 HI[313] NC sky130_fd_sc_hd__conb_1
X\insts[314]  vssd1 vssd1 vccd1 vccd1 HI[314] NC sky130_fd_sc_hd__conb_1
X\insts[315]  vssd1 vssd1 vccd1 vccd1 HI[315] NC sky130_fd_sc_hd__conb_1
X\insts[316]  vssd1 vssd1 vccd1 vccd1 HI[316] NC sky130_fd_sc_hd__conb_1
X\insts[317]  vssd1 vssd1 vccd1 vccd1 HI[317] NC sky130_fd_sc_hd__conb_1
X\insts[318]  vssd1 vssd1 vccd1 vccd1 HI[318] NC sky130_fd_sc_hd__conb_1
X\insts[319]  vssd1 vssd1 vccd1 vccd1 HI[319] NC sky130_fd_sc_hd__conb_1
X\insts[31]  vssd1 vssd1 vccd1 vccd1 HI[31] NC sky130_fd_sc_hd__conb_1
X\insts[320]  vssd1 vssd1 vccd1 vccd1 HI[320] NC sky130_fd_sc_hd__conb_1
X\insts[321]  vssd1 vssd1 vccd1 vccd1 HI[321] NC sky130_fd_sc_hd__conb_1
X\insts[322]  vssd1 vssd1 vccd1 vccd1 HI[322] NC sky130_fd_sc_hd__conb_1
X\insts[323]  vssd1 vssd1 vccd1 vccd1 HI[323] NC sky130_fd_sc_hd__conb_1
X\insts[324]  vssd1 vssd1 vccd1 vccd1 HI[324] NC sky130_fd_sc_hd__conb_1
X\insts[325]  vssd1 vssd1 vccd1 vccd1 HI[325] NC sky130_fd_sc_hd__conb_1
X\insts[326]  vssd1 vssd1 vccd1 vccd1 HI[326] NC sky130_fd_sc_hd__conb_1
X\insts[327]  vssd1 vssd1 vccd1 vccd1 HI[327] NC sky130_fd_sc_hd__conb_1
X\insts[328]  vssd1 vssd1 vccd1 vccd1 HI[328] NC sky130_fd_sc_hd__conb_1
X\insts[329]  vssd1 vssd1 vccd1 vccd1 HI[329] NC sky130_fd_sc_hd__conb_1
X\insts[32]  vssd1 vssd1 vccd1 vccd1 HI[32] NC sky130_fd_sc_hd__conb_1
X\insts[330]  vssd1 vssd1 vccd1 vccd1 HI[330] NC sky130_fd_sc_hd__conb_1
X\insts[331]  vssd1 vssd1 vccd1 vccd1 HI[331] NC sky130_fd_sc_hd__conb_1
X\insts[332]  vssd1 vssd1 vccd1 vccd1 HI[332] NC sky130_fd_sc_hd__conb_1
X\insts[333]  vssd1 vssd1 vccd1 vccd1 HI[333] NC sky130_fd_sc_hd__conb_1
X\insts[334]  vssd1 vssd1 vccd1 vccd1 HI[334] NC sky130_fd_sc_hd__conb_1
X\insts[335]  vssd1 vssd1 vccd1 vccd1 HI[335] NC sky130_fd_sc_hd__conb_1
X\insts[336]  vssd1 vssd1 vccd1 vccd1 HI[336] NC sky130_fd_sc_hd__conb_1
X\insts[337]  vssd1 vssd1 vccd1 vccd1 HI[337] NC sky130_fd_sc_hd__conb_1
X\insts[338]  vssd1 vssd1 vccd1 vccd1 HI[338] NC sky130_fd_sc_hd__conb_1
X\insts[339]  vssd1 vssd1 vccd1 vccd1 HI[339] NC sky130_fd_sc_hd__conb_1
X\insts[33]  vssd1 vssd1 vccd1 vccd1 HI[33] NC sky130_fd_sc_hd__conb_1
X\insts[340]  vssd1 vssd1 vccd1 vccd1 HI[340] NC sky130_fd_sc_hd__conb_1
X\insts[341]  vssd1 vssd1 vccd1 vccd1 HI[341] NC sky130_fd_sc_hd__conb_1
X\insts[342]  vssd1 vssd1 vccd1 vccd1 HI[342] NC sky130_fd_sc_hd__conb_1
X\insts[343]  vssd1 vssd1 vccd1 vccd1 HI[343] NC sky130_fd_sc_hd__conb_1
X\insts[344]  vssd1 vssd1 vccd1 vccd1 HI[344] NC sky130_fd_sc_hd__conb_1
X\insts[345]  vssd1 vssd1 vccd1 vccd1 HI[345] NC sky130_fd_sc_hd__conb_1
X\insts[346]  vssd1 vssd1 vccd1 vccd1 HI[346] NC sky130_fd_sc_hd__conb_1
X\insts[347]  vssd1 vssd1 vccd1 vccd1 HI[347] NC sky130_fd_sc_hd__conb_1
X\insts[348]  vssd1 vssd1 vccd1 vccd1 HI[348] NC sky130_fd_sc_hd__conb_1
X\insts[349]  vssd1 vssd1 vccd1 vccd1 HI[349] NC sky130_fd_sc_hd__conb_1
X\insts[34]  vssd1 vssd1 vccd1 vccd1 HI[34] NC sky130_fd_sc_hd__conb_1
X\insts[350]  vssd1 vssd1 vccd1 vccd1 HI[350] NC sky130_fd_sc_hd__conb_1
X\insts[351]  vssd1 vssd1 vccd1 vccd1 HI[351] NC sky130_fd_sc_hd__conb_1
X\insts[352]  vssd1 vssd1 vccd1 vccd1 HI[352] NC sky130_fd_sc_hd__conb_1
X\insts[353]  vssd1 vssd1 vccd1 vccd1 HI[353] NC sky130_fd_sc_hd__conb_1
X\insts[354]  vssd1 vssd1 vccd1 vccd1 HI[354] NC sky130_fd_sc_hd__conb_1
X\insts[355]  vssd1 vssd1 vccd1 vccd1 HI[355] NC sky130_fd_sc_hd__conb_1
X\insts[356]  vssd1 vssd1 vccd1 vccd1 HI[356] NC sky130_fd_sc_hd__conb_1
X\insts[357]  vssd1 vssd1 vccd1 vccd1 HI[357] NC sky130_fd_sc_hd__conb_1
X\insts[358]  vssd1 vssd1 vccd1 vccd1 HI[358] NC sky130_fd_sc_hd__conb_1
X\insts[359]  vssd1 vssd1 vccd1 vccd1 HI[359] NC sky130_fd_sc_hd__conb_1
X\insts[35]  vssd1 vssd1 vccd1 vccd1 HI[35] NC sky130_fd_sc_hd__conb_1
X\insts[360]  vssd1 vssd1 vccd1 vccd1 HI[360] NC sky130_fd_sc_hd__conb_1
X\insts[361]  vssd1 vssd1 vccd1 vccd1 HI[361] NC sky130_fd_sc_hd__conb_1
X\insts[362]  vssd1 vssd1 vccd1 vccd1 HI[362] NC sky130_fd_sc_hd__conb_1
X\insts[363]  vssd1 vssd1 vccd1 vccd1 HI[363] NC sky130_fd_sc_hd__conb_1
X\insts[364]  vssd1 vssd1 vccd1 vccd1 HI[364] NC sky130_fd_sc_hd__conb_1
X\insts[365]  vssd1 vssd1 vccd1 vccd1 HI[365] NC sky130_fd_sc_hd__conb_1
X\insts[366]  vssd1 vssd1 vccd1 vccd1 HI[366] NC sky130_fd_sc_hd__conb_1
X\insts[367]  vssd1 vssd1 vccd1 vccd1 HI[367] NC sky130_fd_sc_hd__conb_1
X\insts[368]  vssd1 vssd1 vccd1 vccd1 HI[368] NC sky130_fd_sc_hd__conb_1
X\insts[369]  vssd1 vssd1 vccd1 vccd1 HI[369] NC sky130_fd_sc_hd__conb_1
X\insts[36]  vssd1 vssd1 vccd1 vccd1 HI[36] NC sky130_fd_sc_hd__conb_1
X\insts[370]  vssd1 vssd1 vccd1 vccd1 HI[370] NC sky130_fd_sc_hd__conb_1
X\insts[371]  vssd1 vssd1 vccd1 vccd1 HI[371] NC sky130_fd_sc_hd__conb_1
X\insts[372]  vssd1 vssd1 vccd1 vccd1 HI[372] NC sky130_fd_sc_hd__conb_1
X\insts[373]  vssd1 vssd1 vccd1 vccd1 HI[373] NC sky130_fd_sc_hd__conb_1
X\insts[374]  vssd1 vssd1 vccd1 vccd1 HI[374] NC sky130_fd_sc_hd__conb_1
X\insts[375]  vssd1 vssd1 vccd1 vccd1 HI[375] NC sky130_fd_sc_hd__conb_1
X\insts[376]  vssd1 vssd1 vccd1 vccd1 HI[376] NC sky130_fd_sc_hd__conb_1
X\insts[377]  vssd1 vssd1 vccd1 vccd1 HI[377] NC sky130_fd_sc_hd__conb_1
X\insts[378]  vssd1 vssd1 vccd1 vccd1 HI[378] NC sky130_fd_sc_hd__conb_1
X\insts[379]  vssd1 vssd1 vccd1 vccd1 HI[379] NC sky130_fd_sc_hd__conb_1
X\insts[37]  vssd1 vssd1 vccd1 vccd1 HI[37] NC sky130_fd_sc_hd__conb_1
X\insts[380]  vssd1 vssd1 vccd1 vccd1 HI[380] NC sky130_fd_sc_hd__conb_1
X\insts[381]  vssd1 vssd1 vccd1 vccd1 HI[381] NC sky130_fd_sc_hd__conb_1
X\insts[382]  vssd1 vssd1 vccd1 vccd1 HI[382] NC sky130_fd_sc_hd__conb_1
X\insts[383]  vssd1 vssd1 vccd1 vccd1 HI[383] NC sky130_fd_sc_hd__conb_1
X\insts[384]  vssd1 vssd1 vccd1 vccd1 HI[384] NC sky130_fd_sc_hd__conb_1
X\insts[385]  vssd1 vssd1 vccd1 vccd1 HI[385] NC sky130_fd_sc_hd__conb_1
X\insts[386]  vssd1 vssd1 vccd1 vccd1 HI[386] NC sky130_fd_sc_hd__conb_1
X\insts[387]  vssd1 vssd1 vccd1 vccd1 HI[387] NC sky130_fd_sc_hd__conb_1
X\insts[388]  vssd1 vssd1 vccd1 vccd1 HI[388] NC sky130_fd_sc_hd__conb_1
X\insts[389]  vssd1 vssd1 vccd1 vccd1 HI[389] NC sky130_fd_sc_hd__conb_1
X\insts[38]  vssd1 vssd1 vccd1 vccd1 HI[38] NC sky130_fd_sc_hd__conb_1
X\insts[390]  vssd1 vssd1 vccd1 vccd1 HI[390] NC sky130_fd_sc_hd__conb_1
X\insts[391]  vssd1 vssd1 vccd1 vccd1 HI[391] NC sky130_fd_sc_hd__conb_1
X\insts[392]  vssd1 vssd1 vccd1 vccd1 HI[392] NC sky130_fd_sc_hd__conb_1
X\insts[393]  vssd1 vssd1 vccd1 vccd1 HI[393] NC sky130_fd_sc_hd__conb_1
X\insts[394]  vssd1 vssd1 vccd1 vccd1 HI[394] NC sky130_fd_sc_hd__conb_1
X\insts[395]  vssd1 vssd1 vccd1 vccd1 HI[395] NC sky130_fd_sc_hd__conb_1
X\insts[396]  vssd1 vssd1 vccd1 vccd1 HI[396] NC sky130_fd_sc_hd__conb_1
X\insts[397]  vssd1 vssd1 vccd1 vccd1 HI[397] NC sky130_fd_sc_hd__conb_1
X\insts[398]  vssd1 vssd1 vccd1 vccd1 HI[398] NC sky130_fd_sc_hd__conb_1
X\insts[399]  vssd1 vssd1 vccd1 vccd1 HI[399] NC sky130_fd_sc_hd__conb_1
X\insts[39]  vssd1 vssd1 vccd1 vccd1 HI[39] NC sky130_fd_sc_hd__conb_1
X\insts[3]  vssd1 vssd1 vccd1 vccd1 HI[3] NC sky130_fd_sc_hd__conb_1
X\insts[400]  vssd1 vssd1 vccd1 vccd1 HI[400] NC sky130_fd_sc_hd__conb_1
X\insts[401]  vssd1 vssd1 vccd1 vccd1 HI[401] NC sky130_fd_sc_hd__conb_1
X\insts[402]  vssd1 vssd1 vccd1 vccd1 HI[402] NC sky130_fd_sc_hd__conb_1
X\insts[403]  vssd1 vssd1 vccd1 vccd1 HI[403] NC sky130_fd_sc_hd__conb_1
X\insts[404]  vssd1 vssd1 vccd1 vccd1 HI[404] NC sky130_fd_sc_hd__conb_1
X\insts[405]  vssd1 vssd1 vccd1 vccd1 HI[405] NC sky130_fd_sc_hd__conb_1
X\insts[406]  vssd1 vssd1 vccd1 vccd1 HI[406] NC sky130_fd_sc_hd__conb_1
X\insts[407]  vssd1 vssd1 vccd1 vccd1 HI[407] NC sky130_fd_sc_hd__conb_1
X\insts[408]  vssd1 vssd1 vccd1 vccd1 HI[408] NC sky130_fd_sc_hd__conb_1
X\insts[409]  vssd1 vssd1 vccd1 vccd1 HI[409] NC sky130_fd_sc_hd__conb_1
X\insts[40]  vssd1 vssd1 vccd1 vccd1 HI[40] NC sky130_fd_sc_hd__conb_1
X\insts[410]  vssd1 vssd1 vccd1 vccd1 HI[410] NC sky130_fd_sc_hd__conb_1
X\insts[411]  vssd1 vssd1 vccd1 vccd1 HI[411] NC sky130_fd_sc_hd__conb_1
X\insts[412]  vssd1 vssd1 vccd1 vccd1 HI[412] NC sky130_fd_sc_hd__conb_1
X\insts[413]  vssd1 vssd1 vccd1 vccd1 HI[413] NC sky130_fd_sc_hd__conb_1
X\insts[414]  vssd1 vssd1 vccd1 vccd1 HI[414] NC sky130_fd_sc_hd__conb_1
X\insts[415]  vssd1 vssd1 vccd1 vccd1 HI[415] NC sky130_fd_sc_hd__conb_1
X\insts[416]  vssd1 vssd1 vccd1 vccd1 HI[416] NC sky130_fd_sc_hd__conb_1
X\insts[417]  vssd1 vssd1 vccd1 vccd1 HI[417] NC sky130_fd_sc_hd__conb_1
X\insts[418]  vssd1 vssd1 vccd1 vccd1 HI[418] NC sky130_fd_sc_hd__conb_1
X\insts[419]  vssd1 vssd1 vccd1 vccd1 HI[419] NC sky130_fd_sc_hd__conb_1
X\insts[41]  vssd1 vssd1 vccd1 vccd1 HI[41] NC sky130_fd_sc_hd__conb_1
X\insts[420]  vssd1 vssd1 vccd1 vccd1 HI[420] NC sky130_fd_sc_hd__conb_1
X\insts[421]  vssd1 vssd1 vccd1 vccd1 HI[421] NC sky130_fd_sc_hd__conb_1
X\insts[422]  vssd1 vssd1 vccd1 vccd1 HI[422] NC sky130_fd_sc_hd__conb_1
X\insts[423]  vssd1 vssd1 vccd1 vccd1 HI[423] NC sky130_fd_sc_hd__conb_1
X\insts[424]  vssd1 vssd1 vccd1 vccd1 HI[424] NC sky130_fd_sc_hd__conb_1
X\insts[425]  vssd1 vssd1 vccd1 vccd1 HI[425] NC sky130_fd_sc_hd__conb_1
X\insts[426]  vssd1 vssd1 vccd1 vccd1 HI[426] NC sky130_fd_sc_hd__conb_1
X\insts[427]  vssd1 vssd1 vccd1 vccd1 HI[427] NC sky130_fd_sc_hd__conb_1
X\insts[428]  vssd1 vssd1 vccd1 vccd1 HI[428] NC sky130_fd_sc_hd__conb_1
X\insts[429]  vssd1 vssd1 vccd1 vccd1 HI[429] NC sky130_fd_sc_hd__conb_1
X\insts[42]  vssd1 vssd1 vccd1 vccd1 HI[42] NC sky130_fd_sc_hd__conb_1
X\insts[430]  vssd1 vssd1 vccd1 vccd1 HI[430] NC sky130_fd_sc_hd__conb_1
X\insts[431]  vssd1 vssd1 vccd1 vccd1 HI[431] NC sky130_fd_sc_hd__conb_1
X\insts[432]  vssd1 vssd1 vccd1 vccd1 HI[432] NC sky130_fd_sc_hd__conb_1
X\insts[433]  vssd1 vssd1 vccd1 vccd1 HI[433] NC sky130_fd_sc_hd__conb_1
X\insts[434]  vssd1 vssd1 vccd1 vccd1 HI[434] NC sky130_fd_sc_hd__conb_1
X\insts[435]  vssd1 vssd1 vccd1 vccd1 HI[435] NC sky130_fd_sc_hd__conb_1
X\insts[436]  vssd1 vssd1 vccd1 vccd1 HI[436] NC sky130_fd_sc_hd__conb_1
X\insts[437]  vssd1 vssd1 vccd1 vccd1 HI[437] NC sky130_fd_sc_hd__conb_1
X\insts[438]  vssd1 vssd1 vccd1 vccd1 HI[438] NC sky130_fd_sc_hd__conb_1
X\insts[439]  vssd1 vssd1 vccd1 vccd1 HI[439] NC sky130_fd_sc_hd__conb_1
X\insts[43]  vssd1 vssd1 vccd1 vccd1 HI[43] NC sky130_fd_sc_hd__conb_1
X\insts[440]  vssd1 vssd1 vccd1 vccd1 HI[440] NC sky130_fd_sc_hd__conb_1
X\insts[441]  vssd1 vssd1 vccd1 vccd1 HI[441] NC sky130_fd_sc_hd__conb_1
X\insts[442]  vssd1 vssd1 vccd1 vccd1 HI[442] NC sky130_fd_sc_hd__conb_1
X\insts[443]  vssd1 vssd1 vccd1 vccd1 HI[443] NC sky130_fd_sc_hd__conb_1
X\insts[444]  vssd1 vssd1 vccd1 vccd1 HI[444] NC sky130_fd_sc_hd__conb_1
X\insts[445]  vssd1 vssd1 vccd1 vccd1 HI[445] NC sky130_fd_sc_hd__conb_1
X\insts[446]  vssd1 vssd1 vccd1 vccd1 HI[446] NC sky130_fd_sc_hd__conb_1
X\insts[447]  vssd1 vssd1 vccd1 vccd1 HI[447] NC sky130_fd_sc_hd__conb_1
X\insts[448]  vssd1 vssd1 vccd1 vccd1 HI[448] NC sky130_fd_sc_hd__conb_1
X\insts[449]  vssd1 vssd1 vccd1 vccd1 HI[449] NC sky130_fd_sc_hd__conb_1
X\insts[44]  vssd1 vssd1 vccd1 vccd1 HI[44] NC sky130_fd_sc_hd__conb_1
X\insts[450]  vssd1 vssd1 vccd1 vccd1 HI[450] NC sky130_fd_sc_hd__conb_1
X\insts[451]  vssd1 vssd1 vccd1 vccd1 HI[451] NC sky130_fd_sc_hd__conb_1
X\insts[452]  vssd1 vssd1 vccd1 vccd1 HI[452] NC sky130_fd_sc_hd__conb_1
X\insts[453]  vssd1 vssd1 vccd1 vccd1 HI[453] NC sky130_fd_sc_hd__conb_1
X\insts[454]  vssd1 vssd1 vccd1 vccd1 HI[454] NC sky130_fd_sc_hd__conb_1
X\insts[455]  vssd1 vssd1 vccd1 vccd1 HI[455] NC sky130_fd_sc_hd__conb_1
X\insts[456]  vssd1 vssd1 vccd1 vccd1 HI[456] NC sky130_fd_sc_hd__conb_1
X\insts[457]  vssd1 vssd1 vccd1 vccd1 HI[457] NC sky130_fd_sc_hd__conb_1
X\insts[458]  vssd1 vssd1 vccd1 vccd1 HI[458] NC sky130_fd_sc_hd__conb_1
X\insts[459]  vssd1 vssd1 vccd1 vccd1 HI[459] NC sky130_fd_sc_hd__conb_1
X\insts[45]  vssd1 vssd1 vccd1 vccd1 HI[45] NC sky130_fd_sc_hd__conb_1
X\insts[460]  vssd1 vssd1 vccd1 vccd1 HI[460] NC sky130_fd_sc_hd__conb_1
X\insts[461]  vssd1 vssd1 vccd1 vccd1 HI[461] NC sky130_fd_sc_hd__conb_1
X\insts[462]  vssd1 vssd1 vccd1 vccd1 HI[462] NC sky130_fd_sc_hd__conb_1
X\insts[46]  vssd1 vssd1 vccd1 vccd1 HI[46] NC sky130_fd_sc_hd__conb_1
X\insts[47]  vssd1 vssd1 vccd1 vccd1 HI[47] NC sky130_fd_sc_hd__conb_1
X\insts[48]  vssd1 vssd1 vccd1 vccd1 HI[48] NC sky130_fd_sc_hd__conb_1
X\insts[49]  vssd1 vssd1 vccd1 vccd1 HI[49] NC sky130_fd_sc_hd__conb_1
X\insts[4]  vssd1 vssd1 vccd1 vccd1 HI[4] NC sky130_fd_sc_hd__conb_1
X\insts[50]  vssd1 vssd1 vccd1 vccd1 HI[50] NC sky130_fd_sc_hd__conb_1
X\insts[51]  vssd1 vssd1 vccd1 vccd1 HI[51] NC sky130_fd_sc_hd__conb_1
X\insts[52]  vssd1 vssd1 vccd1 vccd1 HI[52] NC sky130_fd_sc_hd__conb_1
X\insts[53]  vssd1 vssd1 vccd1 vccd1 HI[53] NC sky130_fd_sc_hd__conb_1
X\insts[54]  vssd1 vssd1 vccd1 vccd1 HI[54] NC sky130_fd_sc_hd__conb_1
X\insts[55]  vssd1 vssd1 vccd1 vccd1 HI[55] NC sky130_fd_sc_hd__conb_1
X\insts[56]  vssd1 vssd1 vccd1 vccd1 HI[56] NC sky130_fd_sc_hd__conb_1
X\insts[57]  vssd1 vssd1 vccd1 vccd1 HI[57] NC sky130_fd_sc_hd__conb_1
X\insts[58]  vssd1 vssd1 vccd1 vccd1 HI[58] NC sky130_fd_sc_hd__conb_1
X\insts[59]  vssd1 vssd1 vccd1 vccd1 HI[59] NC sky130_fd_sc_hd__conb_1
X\insts[5]  vssd1 vssd1 vccd1 vccd1 HI[5] NC sky130_fd_sc_hd__conb_1
X\insts[60]  vssd1 vssd1 vccd1 vccd1 HI[60] NC sky130_fd_sc_hd__conb_1
X\insts[61]  vssd1 vssd1 vccd1 vccd1 HI[61] NC sky130_fd_sc_hd__conb_1
X\insts[62]  vssd1 vssd1 vccd1 vccd1 HI[62] NC sky130_fd_sc_hd__conb_1
X\insts[63]  vssd1 vssd1 vccd1 vccd1 HI[63] NC sky130_fd_sc_hd__conb_1
X\insts[64]  vssd1 vssd1 vccd1 vccd1 HI[64] NC sky130_fd_sc_hd__conb_1
X\insts[65]  vssd1 vssd1 vccd1 vccd1 HI[65] NC sky130_fd_sc_hd__conb_1
X\insts[66]  vssd1 vssd1 vccd1 vccd1 HI[66] NC sky130_fd_sc_hd__conb_1
X\insts[67]  vssd1 vssd1 vccd1 vccd1 HI[67] NC sky130_fd_sc_hd__conb_1
X\insts[68]  vssd1 vssd1 vccd1 vccd1 HI[68] NC sky130_fd_sc_hd__conb_1
X\insts[69]  vssd1 vssd1 vccd1 vccd1 HI[69] NC sky130_fd_sc_hd__conb_1
X\insts[6]  vssd1 vssd1 vccd1 vccd1 HI[6] NC sky130_fd_sc_hd__conb_1
X\insts[70]  vssd1 vssd1 vccd1 vccd1 HI[70] NC sky130_fd_sc_hd__conb_1
X\insts[71]  vssd1 vssd1 vccd1 vccd1 HI[71] NC sky130_fd_sc_hd__conb_1
X\insts[72]  vssd1 vssd1 vccd1 vccd1 HI[72] NC sky130_fd_sc_hd__conb_1
X\insts[73]  vssd1 vssd1 vccd1 vccd1 HI[73] NC sky130_fd_sc_hd__conb_1
X\insts[74]  vssd1 vssd1 vccd1 vccd1 HI[74] NC sky130_fd_sc_hd__conb_1
X\insts[75]  vssd1 vssd1 vccd1 vccd1 HI[75] NC sky130_fd_sc_hd__conb_1
X\insts[76]  vssd1 vssd1 vccd1 vccd1 HI[76] NC sky130_fd_sc_hd__conb_1
X\insts[77]  vssd1 vssd1 vccd1 vccd1 HI[77] NC sky130_fd_sc_hd__conb_1
X\insts[78]  vssd1 vssd1 vccd1 vccd1 HI[78] NC sky130_fd_sc_hd__conb_1
X\insts[79]  vssd1 vssd1 vccd1 vccd1 HI[79] NC sky130_fd_sc_hd__conb_1
X\insts[7]  vssd1 vssd1 vccd1 vccd1 HI[7] NC sky130_fd_sc_hd__conb_1
X\insts[80]  vssd1 vssd1 vccd1 vccd1 HI[80] NC sky130_fd_sc_hd__conb_1
X\insts[81]  vssd1 vssd1 vccd1 vccd1 HI[81] NC sky130_fd_sc_hd__conb_1
X\insts[82]  vssd1 vssd1 vccd1 vccd1 HI[82] NC sky130_fd_sc_hd__conb_1
X\insts[83]  vssd1 vssd1 vccd1 vccd1 HI[83] NC sky130_fd_sc_hd__conb_1
X\insts[84]  vssd1 vssd1 vccd1 vccd1 HI[84] NC sky130_fd_sc_hd__conb_1
X\insts[85]  vssd1 vssd1 vccd1 vccd1 HI[85] NC sky130_fd_sc_hd__conb_1
X\insts[86]  vssd1 vssd1 vccd1 vccd1 HI[86] NC sky130_fd_sc_hd__conb_1
X\insts[87]  vssd1 vssd1 vccd1 vccd1 HI[87] NC sky130_fd_sc_hd__conb_1
X\insts[88]  vssd1 vssd1 vccd1 vccd1 HI[88] NC sky130_fd_sc_hd__conb_1
X\insts[89]  vssd1 vssd1 vccd1 vccd1 HI[89] NC sky130_fd_sc_hd__conb_1
X\insts[8]  vssd1 vssd1 vccd1 vccd1 HI[8] NC sky130_fd_sc_hd__conb_1
X\insts[90]  vssd1 vssd1 vccd1 vccd1 HI[90] NC sky130_fd_sc_hd__conb_1
X\insts[91]  vssd1 vssd1 vccd1 vccd1 HI[91] NC sky130_fd_sc_hd__conb_1
X\insts[92]  vssd1 vssd1 vccd1 vccd1 HI[92] NC sky130_fd_sc_hd__conb_1
X\insts[93]  vssd1 vssd1 vccd1 vccd1 HI[93] NC sky130_fd_sc_hd__conb_1
X\insts[94]  vssd1 vssd1 vccd1 vccd1 HI[94] NC sky130_fd_sc_hd__conb_1
X\insts[95]  vssd1 vssd1 vccd1 vccd1 HI[95] NC sky130_fd_sc_hd__conb_1
X\insts[96]  vssd1 vssd1 vccd1 vccd1 HI[96] NC sky130_fd_sc_hd__conb_1
X\insts[97]  vssd1 vssd1 vccd1 vccd1 HI[97] NC sky130_fd_sc_hd__conb_1
X\insts[98]  vssd1 vssd1 vccd1 vccd1 HI[98] NC sky130_fd_sc_hd__conb_1
X\insts[99]  vssd1 vssd1 vccd1 vccd1 HI[99] NC sky130_fd_sc_hd__conb_1
X\insts[9]  vssd1 vssd1 vccd1 vccd1 HI[9] NC sky130_fd_sc_hd__conb_1

.ends
.end
