* Extracted by KLayout on : 19/01/2022 09:20

.SUBCKT spare_logic_block spare_xz[15] spare_xz[23] spare_xz[26] spare_xz[6]
+ spare_xz[19] spare_xi[1] spare_xno[0] spare_xz[24] spare_xz[16] vccd
+ spare_xz[1] spare_xz[8] spare_xna[1] spare_xz[22] spare_xfqn[1] spare_xfq[1]
+ spare_xz[20] spare_xfq[0] spare_xi[0] spare_xz[21] spare_xz[25] spare_xz[0]
+ spare_xfqn[0] spare_xz[7] spare_xmx[1] spare_xz[9] spare_xz[14] spare_xz[11]
+ spare_xz[18] spare_xz[12] spare_xz[17] spare_xi[3] spare_xz[13] spare_xi[2]
+ spare_xmx[0] spare_xno[1] spare_xz[10] spare_xz[5] spare_xz[3] spare_xz[4]
+ spare_xna[0] spare_xz[2] spare_xib vssd
X$1 vssd spare_xmx[0] spare_xz[13] spare_xz[15] spare_xz[17] vccd vccd vssd
+ sky130_fd_sc_hd__mux2_2
X$2 vccd vccd vssd spare_xz[15] vssd sky130_fd_sc_hd__conb_1
X$3 vssd spare_xz[23] spare_xfqn[0] spare_xfq[0] spare_xz[21] spare_xz[19]
+ spare_xz[25] vccd vccd vssd sky130_fd_sc_hd__dfbbp_1
X$4 vccd vccd vssd spare_xz[23] vssd sky130_fd_sc_hd__conb_1
X$5 vssd spare_xz[24] spare_xfqn[1] spare_xfq[1] spare_xz[22] spare_xz[20]
+ spare_xz[26] vccd vccd vssd sky130_fd_sc_hd__dfbbp_1
X$6 vccd vccd vssd spare_xz[26] vssd sky130_fd_sc_hd__conb_1
X$7 vccd vccd spare_xna[1] spare_xz[8] vssd spare_xz[6] vssd
+ sky130_fd_sc_hd__nand2_2
X$8 vccd vccd vssd spare_xz[6] vssd sky130_fd_sc_hd__conb_1
X$9 vccd vccd vssd spare_xz[19] vssd sky130_fd_sc_hd__conb_1
X$10 vccd vssd vccd spare_xi[1] spare_xz[1] vssd sky130_fd_sc_hd__inv_2
X$11 vccd vssd spare_xz[9] vccd spare_xno[0] spare_xz[11] vssd
+ sky130_fd_sc_hd__nor2_2
X$12 vccd vccd vssd spare_xz[24] vssd sky130_fd_sc_hd__conb_1
X$13 vssd spare_xmx[1] spare_xz[14] spare_xz[16] spare_xz[18] vccd vccd vssd
+ sky130_fd_sc_hd__mux2_2
X$14 vccd vccd vssd spare_xz[16] vssd sky130_fd_sc_hd__conb_1
X$15 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$16 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$17 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$18 vccd vccd vssd spare_xz[21] vssd sky130_fd_sc_hd__conb_1
X$19 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$20 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$21 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$22 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$23 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$24 vccd vccd vssd spare_xz[25] vssd sky130_fd_sc_hd__conb_1
X$25 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$26 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$27 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$28 vccd vssd vccd spare_xi[0] spare_xz[0] vssd sky130_fd_sc_hd__inv_2
X$29 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$30 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$31 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$32 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$33 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$34 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$35 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$36 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$37 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$38 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$39 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$40 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$41 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$42 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$43 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$44 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$45 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$46 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$47 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$48 vccd vccd vssd spare_xz[8] vssd sky130_fd_sc_hd__conb_1
X$49 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$50 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$51 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$52 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$53 vccd vccd vssd spare_xz[1] vssd sky130_fd_sc_hd__conb_1
X$54 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$55 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$56 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$57 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$58 vccd vccd vssd spare_xz[22] vssd sky130_fd_sc_hd__conb_1
X$59 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$60 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$61 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$62 vccd vccd vssd spare_xz[20] vssd sky130_fd_sc_hd__conb_1
X$63 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$64 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$65 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$66 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$67 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$68 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$69 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$70 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$71 vccd vssd spare_xz[10] vccd spare_xno[1] spare_xz[12] vssd
+ sky130_fd_sc_hd__nor2_2
X$72 vccd vccd vssd spare_xz[12] vssd sky130_fd_sc_hd__conb_1
X$73 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$74 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$75 vccd vccd vssd spare_xz[10] vssd sky130_fd_sc_hd__conb_1
X$76 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$77 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$78 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$79 vccd vccd vssd spare_xz[5] vssd sky130_fd_sc_hd__conb_1
X$80 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$81 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$82 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$83 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$84 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$85 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$86 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$87 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$88 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$89 vccd vccd vssd spare_xz[3] vssd sky130_fd_sc_hd__conb_1
X$90 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$91 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$92 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$93 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$94 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$95 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$96 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$97 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$98 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$99 vssd spare_xz[4] spare_xib vccd vccd vssd sky130_fd_sc_hd__inv_8
X$100 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$101 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$102 vccd vccd vssd spare_xz[4] vssd sky130_fd_sc_hd__conb_1
X$103 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$104 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$105 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$106 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$107 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$108 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$109 vccd vccd spare_xna[0] spare_xz[7] vssd spare_xz[5] vssd
+ sky130_fd_sc_hd__nand2_2
X$110 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$111 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$112 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$113 vccd vssd vccd spare_xi[3] spare_xz[3] vssd sky130_fd_sc_hd__inv_2
X$114 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$115 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$116 vccd vccd vssd spare_xz[2] vssd sky130_fd_sc_hd__conb_1
X$117 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$118 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$119 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$120 vccd vccd vssd spare_xz[13] vssd sky130_fd_sc_hd__conb_1
X$121 vccd vssd vccd spare_xi[2] spare_xz[2] vssd sky130_fd_sc_hd__inv_2
X$122 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$123 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$124 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$125 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$126 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$127 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$128 vccd vssd vccd vssd sky130_fd_sc_hd__fill_2
X$129 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$130 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$131 vccd vccd vssd spare_xz[7] vssd sky130_fd_sc_hd__conb_1
X$132 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$133 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$134 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$135 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$136 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$137 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$138 vccd vccd vssd vssd sky130_fd_sc_hd__decap_6
X$139 vccd vccd vssd spare_xz[9] vssd sky130_fd_sc_hd__conb_1
X$140 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$141 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$142 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$143 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$144 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$145 vccd vccd vssd spare_xz[0] vssd sky130_fd_sc_hd__conb_1
X$146 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$147 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$148 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$149 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$150 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$151 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$152 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$153 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$154 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$155 vccd vccd vssd spare_xz[14] vssd sky130_fd_sc_hd__conb_1
X$156 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$157 vccd vccd vssd spare_xz[18] vssd sky130_fd_sc_hd__conb_1
X$158 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$159 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$160 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$161 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$162 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$163 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$164 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$165 vccd vccd vssd vssd sky130_fd_sc_hd__decap_12
X$166 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$167 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$168 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$169 vccd vccd vssd spare_xz[17] vssd sky130_fd_sc_hd__conb_1
X$170 vccd vssd sky130_fd_sc_hd__tapvpwrvgnd_1
X$171 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$172 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$173 vccd vccd vssd vssd sky130_fd_sc_hd__decap_8
X$174 vccd vccd vssd spare_xz[11] vssd sky130_fd_sc_hd__conb_1
X$175 vccd vssd vccd vssd sky130_fd_sc_hd__decap_4
X$176 vccd vssd vccd vssd sky130_fd_sc_hd__fill_1
X$177 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
X$178 vccd vssd vccd vssd sky130_fd_sc_hd__decap_3
.ENDS spare_logic_block

.SUBCKT sky130_fd_sc_hd__nand2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__inv_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_8

.SUBCKT sky130_fd_sc_hd__fill_2 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__inv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__fill_1 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__nor2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_2

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 nc_1 nc_2
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__decap_6 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__mux2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_2

.SUBCKT sky130_fd_sc_hd__conb_1 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__decap_3 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__decap_4 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__decap_12 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__decap_8 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__dfbbp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__dfbbp_1
