* Extracted by KLayout on : 19/01/2022 09:20

.SUBCKT gpio_defaults_block gpio_defaults[2] gpio_defaults[4] gpio_defaults[11]
+ VPWR gpio_defaults[1] gpio_defaults[3] gpio_defaults[5] gpio_defaults[9]
+ gpio_defaults[10] gpio_defaults[0] gpio_defaults[6] gpio_defaults[7]
+ gpio_defaults[8] gpio_defaults[12] VGND
X$1 VPWR VPWR VGND gpio_defaults[2] \$I143 VGND sky130_fd_sc_hd__conb_1
X$2 VPWR VPWR VGND gpio_defaults[4] \$I145 VGND sky130_fd_sc_hd__conb_1
X$3 VPWR VPWR VGND gpio_defaults[11] \$I137 VGND sky130_fd_sc_hd__conb_1
X$4 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$5 VPWR VPWR VGND gpio_defaults[7] \$I136 VGND sky130_fd_sc_hd__conb_1
X$6 VPWR VPWR VGND gpio_defaults[8] \$I140 VGND sky130_fd_sc_hd__conb_1
X$7 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$8 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$9 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$10 VPWR VPWR VGND gpio_defaults[6] \$I142 VGND sky130_fd_sc_hd__conb_1
X$11 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$12 VPWR VPWR VGND gpio_defaults[9] \$I141 VGND sky130_fd_sc_hd__conb_1
X$13 VPWR VPWR VGND gpio_defaults[5] \$I146 VGND sky130_fd_sc_hd__conb_1
X$14 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$15 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$16 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$17 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$18 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$19 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$20 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$21 VPWR VPWR VGND gpio_defaults[0] \$I147 VGND sky130_fd_sc_hd__conb_1
X$22 VPWR VPWR VGND \$I133 gpio_defaults[1] VGND sky130_fd_sc_hd__conb_1
X$23 VPWR VPWR VGND gpio_defaults[3] \$I144 VGND sky130_fd_sc_hd__conb_1
X$24 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$25 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$26 VPWR VPWR VGND gpio_defaults[12] \$I139 VGND sky130_fd_sc_hd__conb_1
X$27 VPWR VPWR VGND \$I126 gpio_defaults[10] VGND sky130_fd_sc_hd__conb_1
X$28 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$29 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$30 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$31 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_2
X$32 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$33 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$34 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$35 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$36 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$37 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$38 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$39 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$40 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
X$41 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$42 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$43 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$44 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$45 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$46 VPWR VGND VPWR VGND sky130_fd_sc_hd__fill_1
X$47 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$48 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$49 VPWR VGND sky130_fd_sc_hd__tapvpwrvgnd_1
.ENDS gpio_defaults_block

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 nc_1 nc_2
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__decap_3 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__decap_4 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__fill_1 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__decap_12 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__conb_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__fill_2 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__decap_6 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_6
