*
*  /home/marwan/ef/klayout_lvs/lvs/test_cases/mprj_logic_high/mprj_logic_high.spice : SPICE netlist translated from the VERILOG netlist : /home/marwan/ef/caravel/verilog/gl/mprj_logic_high.v
*                                                                                     on the 2021-12-22 17:57:47.045915
*
************************************************************************************************************************************************************************************************

.INCLUDE sky130_fd_sc_hd.spice 

.GLOBAL VDD VSS

.SUBCKT MPRJ_LOGIC_HIGH VCCD1 VSSD1 HI[0] HI[1] HI[2] HI[3] HI[4] HI[5] HI[6] HI[7] HI[8] HI[9] HI[10] HI[11] HI[12] HI[13] HI[14] HI[15] HI[16] HI[17] HI[18] HI[19] HI[20] HI[21] HI[22] HI[23] HI[24] HI[25] HI[26] HI[27] HI[28] HI[29] HI[30] HI[31] HI[32] HI[33] HI[34] HI[35] HI[36] HI[37] HI[38] HI[39] HI[40] HI[41] HI[42] HI[43] HI[44] HI[45] HI[46] HI[47] HI[48] HI[49] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58] HI[59] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[90] HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106] HI[107] HI[108] HI[109] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116] HI[117] HI[118] HI[119] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126] HI[127] HI[128] HI[129] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136] HI[137] HI[138] HI[139] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146] HI[147] HI[148] HI[149] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156] HI[157] HI[158] HI[159] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166] HI[167] HI[168] HI[169] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176] HI[177] HI[178] HI[179] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186] HI[187] HI[188] HI[189] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196] HI[197] HI[198] HI[199] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205] HI[206] HI[207] HI[208] HI[209] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215] HI[216] HI[217] HI[218] HI[219] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225] HI[226] HI[227] HI[228] HI[229] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235] HI[236] HI[237] HI[238] HI[239] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245] HI[246] HI[247] HI[248] HI[249] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255] HI[256] HI[257] HI[258] HI[259] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265] HI[266] HI[267] HI[268] HI[269] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275] HI[276] HI[277] HI[278] HI[279] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285] HI[286] HI[287] HI[288] HI[289] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295] HI[296] HI[297] HI[298] HI[299] HI[300] HI[301] HI[302] HI[303] HI[304] HI[305] HI[306] HI[307] HI[308] HI[309] HI[310] HI[311] HI[312] HI[313] HI[314] HI[315] HI[316] HI[317] HI[318] HI[319] HI[320] HI[321] HI[322] HI[323] HI[324] HI[325] HI[326] HI[327] HI[328] HI[329] HI[330] HI[331] HI[332] HI[333] HI[334] HI[335] HI[336] HI[337] HI[338] HI[339] HI[340] HI[341] HI[342] HI[343] HI[344] HI[345] HI[346] HI[347] HI[348] HI[349] HI[350] HI[351] HI[352] HI[353] HI[354] HI[355] HI[356] HI[357] HI[358] HI[359] HI[360] HI[361] HI[362] HI[363] HI[364] HI[365] HI[366] HI[367] HI[368] HI[369] HI[370] HI[371] HI[372] HI[373] HI[374] HI[375] HI[376] HI[377] HI[378] HI[379] HI[380] HI[381] HI[382] HI[383] HI[384] HI[385] HI[386] HI[387] HI[388] HI[389] HI[390] HI[391] HI[392] HI[393] HI[394] HI[395] HI[396] HI[397] HI[398] HI[399] HI[400] HI[401] HI[402] HI[403] HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[410] HI[411] HI[412] HI[413] HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[420] HI[421] HI[422] HI[423] HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[430] HI[431] HI[432] HI[433] HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[440] HI[441] HI[442] HI[443] HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[450] HI[451] HI[452] HI[453] HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[460] HI[461] HI[462] 

XFILLER_0_111 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_119 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_139 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_141 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_166 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_172 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_194 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_228 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_245 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_259 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_279 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_284 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_29 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_3 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_306 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_309 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_334 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_421 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_446 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_458 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_474 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_483 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_502 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_55 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_57 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_601 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_613 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_0_617 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_629 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_641 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_0_645 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_657 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_669 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_0_67 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_673 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_685 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_697 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_0_701 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_713 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_0_725 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_0_729 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_0_77 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_0_94 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_108 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_1_113 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_1_117 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_121 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_133 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_142 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_154 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_166 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_172 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_184 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_196 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_1_204 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_209 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_221 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_1_225 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_230 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_242 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_254 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_1_261 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_273 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_279 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_281 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_293 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_1_3 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_1_301 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_1_307 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_319 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_1_327 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_331 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_1_335 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_337 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_1_343 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_355 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_367 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_379 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_391 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_393 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_405 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_417 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_429 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_441 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_447 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_449 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_461 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_467 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_471 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_1_479 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_484 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_1_490 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_502 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_505 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_517 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_529 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_541 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_55 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_553 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_557 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_1_561 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_573 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_585 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_597 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_609 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_615 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_617 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_629 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_63 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_641 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_653 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_665 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_671 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_673 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_68 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_685 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_697 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_709 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_721 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_1_727 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_729 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_1_80 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_1_92 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_1_96 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_109 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_11 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_118 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_130 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_138 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_141 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_153 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_165 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_177 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_189 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_195 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_197 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_209 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_221 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_233 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_245 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_251 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_253 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_265 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_277 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_289 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_29 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_297 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_3 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_302 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_309 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_321 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_333 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_345 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_357 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_363 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_365 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_377 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_386 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_398 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_410 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_418 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_421 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_433 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_442 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_454 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_466 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_470 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_477 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_502 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_514 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_52 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_526 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_533 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_545 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_557 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_569 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_581 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_587 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_589 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_60 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_601 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_613 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_625 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_637 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_2_643 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_645 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_657 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_669 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_681 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_689 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XFILLER_2_695 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_2_710 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_72 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_722 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_8
XFILLER_2_730 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_2_85 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_2_97 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_3_116 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_139 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_3_141 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_3_166 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_29 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_3 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_3_40 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_3_486 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_12
XFILLER_3_498 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_3_50 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XFILLER_3_511 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_4
XFILLER_3_530 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_54 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_722 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_6
XFILLER_3_729 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_2
XFILLER_3_9 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__FILL_1
XPHY_0 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_1 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_2 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_3 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_4 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_5 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_6 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XPHY_7 VSSD1 VSSD1 VCCD1 VCCD1 SKY130_FD_SC_HD__DECAP_3
XTAP_10 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_11 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_12 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_13 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_14 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_15 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_16 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_17 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_18 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_19 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_20 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_21 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_22 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_23 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_24 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_25 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_26 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_27 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_28 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_29 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_30 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_31 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_32 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_33 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_34 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_35 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_36 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_37 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_38 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_39 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_40 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_41 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_42 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_43 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_44 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_45 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_46 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_47 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_48 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_49 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_50 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_51 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_52 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_53 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_54 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_55 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_56 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_57 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_58 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_59 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_60 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_61 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_62 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_63 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_64 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_65 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_66 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_67 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_68 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_69 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_70 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_71 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_72 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_73 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_74 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_75 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_76 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_77 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_78 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_79 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_8 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_80 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_81 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_82 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_83 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_84 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_85 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_9 VSSD1 VCCD1 SKY130_FD_SC_HD__TAPVPWRVGND_1
