*
*  /home/marwan/KLayout_Support_for_Sky130A/LVS/test_cases/digital_pll/digital_pll.spice : SPICE netlist translated from the VERILOG netlist : /home/marwan/caravel/verilog/gl/digital_pll.v
*                                                                                          on the 2021-12-20 06:29:16.007670
*
**********************************************************************************************************************************************************************************************

.INCLUDE sky130_fd_sc_hd_new.spice 

.GLOBAL VDD VSS

.SUBCKT DIGITAL_PLL VGND VPWR DCO ENABLE OSC RESETB CLOCKP[0] CLOCKP[1] DIV[0] DIV[1] DIV[2] DIV[3] DIV[4] EXT_TRIM[0] EXT_TRIM[1] EXT_TRIM[2] EXT_TRIM[3] EXT_TRIM[4] EXT_TRIM[5] EXT_TRIM[6] EXT_TRIM[7] EXT_TRIM[8] EXT_TRIM[9] EXT_TRIM[10] EXT_TRIM[11] EXT_TRIM[12] EXT_TRIM[13] EXT_TRIM[14] EXT_TRIM[15] EXT_TRIM[16] EXT_TRIM[17] EXT_TRIM[18] EXT_TRIM[19] EXT_TRIM[20] EXT_TRIM[21] EXT_TRIM[22] EXT_TRIM[23] EXT_TRIM[24] EXT_TRIM[25] 

XANTENNA__177__A DIV[0] VGND VNB VPB VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__181__A ENABLE VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__181__B RESETB VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__182__A DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__201__A1 DIV[3] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__201__B1 DIV[2] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__202__A DIV[3] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__204__A1 DIV[2] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__207__A DIV[1] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__210__A1 DIV[1] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__210__B1 DIV[0] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__211__A1 DIV[1] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__216__A DIV[4] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__218__B1 DIV[4] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__330__A1 EXT_TRIM[11] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__330__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__331__A1 EXT_TRIM[24] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__331__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__332__A1 EXT_TRIM[10] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__332__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__333__A1 EXT_TRIM[23] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__333__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__334__A1 EXT_TRIM[9] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__334__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__335__A1 EXT_TRIM[22] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__335__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__336__A1 EXT_TRIM[8] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__336__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__337__A1 EXT_TRIM[21] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__337__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__338__A1 EXT_TRIM[7] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__338__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__339__A1 EXT_TRIM[20] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__339__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__340__A1 EXT_TRIM[6] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__340__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__341__A1 EXT_TRIM[19] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__341__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__342__A1 EXT_TRIM[5] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__342__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__343__A1 EXT_TRIM[18] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__343__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__344__A1 EXT_TRIM[4] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__344__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__345__A1 EXT_TRIM[17] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__345__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__346__A1 EXT_TRIM[3] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__346__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__347__A1 EXT_TRIM[16] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__347__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__348__A1 EXT_TRIM[2] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__348__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__349__A1 EXT_TRIM[15] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__349__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__350__A1 EXT_TRIM[1] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__350__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__351__A1 EXT_TRIM[14] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__351__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__352__A1 EXT_TRIM[0] VPWR VGND VPWR VGND SKY130_FD_SC_HD__DIODE_2
XANTENNA__352__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__353__A1 EXT_TRIM[13] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__353__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__354__A1 EXT_TRIM[12] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__354__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__355__A1 EXT_TRIM[25] VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__355__S DCO VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XANTENNA__356__D OSC VGND VGND VPWR VPWR SKY130_FD_SC_HD__DIODE_2
XFILLER_0_10 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_0_105 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_0_19 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_0_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_0_37 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_0_52 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_0_62 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_0_66 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_0_70 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_0_82 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_0_93 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_10_10 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_10_104 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_10_19 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_10_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_10_36 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_10_7 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_10_94 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_11_101 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_11_111 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_11_130 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_11_23 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_11_32 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_11_38 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_11_50 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_11_57 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_11_77 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_12_101 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_12_105 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_12_19 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_12_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_12_39 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_12_48 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_12_68 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_12_80 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_13_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_13_34 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_13_54 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_14_112 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_14_13 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_14_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_14_43 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_14_63 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_14_81 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_14_85 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_15_109 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_15_24 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_15_39 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_15_5 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_15_53 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_15_67 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_15_76 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_15_93 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_8
XFILLER_16_115 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_16_135 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_16_23 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_16_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_16_32 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_16_59 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_16_7 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_16_72 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_16_94 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_16_98 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_17_100 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_17_12 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_17_30 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_18_112 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_18_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_18_26 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_18_49 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_18_75 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_18_96 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_100 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_120 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_135 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_28 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_55 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_68 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_19_87 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_1_111 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_1_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_1_54 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_1_78 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_20_112 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_20_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_20_38 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_20_5 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_21_104 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_21_135 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_21_21 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_21_55 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_21_69 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_22_133 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_22_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_22_31 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_22_42 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_22_7 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_22_72 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_2_120 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_2_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_2_18 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_2_5 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_2_78 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_3_111 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_3_113 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_3_28 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_3_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_3_33 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_3_37 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_3_48 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_3_57 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_3_71 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_3_94 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_4_120 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_4_129 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_4_135 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_4_58 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_4_81 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_5_103 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_5_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_5_19 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_5_32 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_5_57 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_5_69 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_6_100 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_6_122 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_6_134 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_6_17 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_6_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_6_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_6_38 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_6_53 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_6_62 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_4
XFILLER_6_71 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_6_83 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_6_88 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_7_103 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_7_116 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_8
XFILLER_7_127 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_8
XFILLER_7_135 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_7_39 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XFILLER_7_81 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_7_90 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_7_96 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_8_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_8_29 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_8_51 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_12
XFILLER_8_63 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_6
XFILLER_8_69 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_9_113 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_9_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_9_47 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_2
XFILLER_9_5 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_9_52 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_9_78 VGND VGND VPWR VPWR SKY130_FD_SC_HD__FILL_1
XFILLER_9_87 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_0 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_1 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_10 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_11 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_12 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_13 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_14 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_15 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_16 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_17 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_18 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_19 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_2 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_20 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_21 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_22 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_23 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_24 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_25 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_26 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_27 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_28 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_29 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_3 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_30 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_31 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_32 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_33 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_34 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_35 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_36 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_37 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_38 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_39 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_4 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_40 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_41 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_42 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_43 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_44 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_45 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_5 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_6 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_7 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_8 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XPHY_9 VGND VGND VPWR VPWR SKY130_FD_SC_HD__DECAP_3
XTAP_46 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_47 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_48 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_49 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_50 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_51 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_52 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_53 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_54 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_55 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_56 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_57 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_58 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_59 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_60 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_61 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_62 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_63 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_64 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_65 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_66 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_67 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_68 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_69 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_70 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_71 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_72 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_73 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_74 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_75 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_76 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_77 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_78 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_79 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_80 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_81 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_82 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_83 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_84 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_85 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_86 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_87 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_88 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_89 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_90 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_91 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_92 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_93 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_94 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
XTAP_95 VGND VPWR SKY130_FD_SC_HD__TAPVPWRVGND_1
X_164_ \PLL_CONTRO VGND VGND VPWR VPWR _072_ SKY130_FD_SC_HD__INV_2
X_165_ \PLL_CONTRO VGND VGND VPWR VPWR _073_ SKY130_FD_SC_HD__INV_2
X_166_ \PLL_CONTRO VGND VGND VPWR VPWR _074_ SKY130_FD_SC_HD__INV_2
X_167_ \PLL_CONTRO VGND VGND VPWR VPWR _075_ SKY130_FD_SC_HD__INV_2
X_168_ \PLL_CONTRO VGND VGND VPWR VPWR _076_ SKY130_FD_SC_HD__INV_2
X_169_ \PLL_CONTRO VGND VGND VPWR VPWR _077_ SKY130_FD_SC_HD__INV_2
X_170_ \PLL_CONTRO VGND VGND VPWR VPWR _078_ SKY130_FD_SC_HD__INV_2
X_171_ \PLL_CONTRO VGND VGND VPWR VPWR _079_ SKY130_FD_SC_HD__INV_2
X_172_ \PLL_CONTRO VGND VGND VPWR VPWR _080_ SKY130_FD_SC_HD__INV_2
X_173_ \PLL_CONTRO VGND VGND VPWR VPWR _081_ SKY130_FD_SC_HD__INV_2
X_174_ \PLL_CONTRO VGND VGND VPWR VPWR _082_ SKY130_FD_SC_HD__INV_2
X_175_ \PLL_CONTRO VGND VGND VPWR VPWR _083_ SKY130_FD_SC_HD__INV_2
X_176_ \PLL_CONTRO VGND VGND VPWR VPWR _084_ SKY130_FD_SC_HD__INV_2
X_177_ DIV[0] VGND VGND VPWR VPWR _085_ SKY130_FD_SC_HD__INV_2
X_178_ \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _086_ SKY130_FD_SC_HD__A2BB2O_2
X_179_ _086_ VGND VGND VPWR VPWR _087_ SKY130_FD_SC_HD__INV_2
X_180_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _071_ SKY130_FD_SC_HD__A22O_2
X_181_ ENABLE RESETB VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__NAND2_2
X_182_ DCO \RINGOS VGND VGND VPWR VPWR _050_ SKY130_FD_SC_HD__NOR2_2
X_183_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _070_ SKY130_FD_SC_HD__A22O_2
X_184_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _069_ SKY130_FD_SC_HD__A22O_2
X_185_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _068_ SKY130_FD_SC_HD__A22O_2
X_186_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _067_ SKY130_FD_SC_HD__A22O_2
X_187_ \PLL_CONTRO _087_ \PLL_CONTRO _086_ VGND VGND VPWR VPWR _066_ SKY130_FD_SC_HD__A22O_2
X_188_ \PLL_CONTRO _086_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _065_ SKY130_FD_SC_HD__A22O_2
X_189_ \PLL_CONTRO _087_ VGND VGND VPWR VPWR _064_ SKY130_FD_SC_HD__OR2_2
X_190_ \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _088_ SKY130_FD_SC_HD__NOR2_2
X_191_ \PLL_CONTRO \PLL_CONTRO _088_ VGND VGND VPWR VPWR _089_ SKY130_FD_SC_HD__A21O_2
X_192_ \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _090_ SKY130_FD_SC_HD__NOR2_2
X_193_ _076_ _077_ VGND VGND VPWR VPWR _091_ SKY130_FD_SC_HD__NOR2_2
X_194_ \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _092_ SKY130_FD_SC_HD__O2BB2A_2
X_195_ \PLL_CONTRO \PLL_CONTRO _091_ _092_ VGND VGND VPWR VPWR _093_ SKY130_FD_SC_HD__A22O_2
X_196_ _093_ VGND VGND VPWR VPWR _094_ SKY130_FD_SC_HD__INV_2
X_197_ \PLL_CONTRO \PLL_CONTRO _090_ _094_ VGND VGND VPWR VPWR _095_ SKY130_FD_SC_HD__O2BB2A_2
X_198_ _089_ _095_ _089_ _095_ VGND VGND VPWR VPWR _096_ SKY130_FD_SC_HD__A2BB2O_2
X_199_ \PLL_CONTRO \PLL_CONTRO _090_ VGND VGND VPWR VPWR _097_ SKY130_FD_SC_HD__A21OI_2
X_200_ _093_ _097_ _093_ _097_ VGND VGND VPWR VPWR _098_ SKY130_FD_SC_HD__A2BB2O_2
X_201_ DIV[3] _096_ DIV[2] _098_ VGND VGND VPWR VPWR _099_ SKY130_FD_SC_HD__A22OI_2
X_202_ DIV[3] _096_ VGND VGND VPWR VPWR _100_ SKY130_FD_SC_HD__OR2_2
X_203_ _100_ VGND VGND VPWR VPWR _101_ SKY130_FD_SC_HD__INV_2
X_204_ DIV[2] _098_ _100_ _099_ VGND VGND VPWR VPWR _102_ SKY130_FD_SC_HD__O211A_2
X_205_ _102_ VGND VGND VPWR VPWR _103_ SKY130_FD_SC_HD__INV_2
X_206_ _091_ _092_ _091_ _092_ VGND VGND VPWR VPWR _104_ SKY130_FD_SC_HD__O2BB2AI_2
X_207_ DIV[1] _104_ VGND VGND VPWR VPWR _105_ SKY130_FD_SC_HD__NAND2_2
X_208_ _076_ _077_ _091_ VGND VGND VPWR VPWR _106_ SKY130_FD_SC_HD__A21OI_2
X_209_ _106_ VGND VGND VPWR VPWR _107_ SKY130_FD_SC_HD__INV_2
X_210_ DIV[1] _104_ DIV[0] _107_ _105_ VGND VGND VPWR VPWR _108_ SKY130_FD_SC_HD__O221A_2
X_211_ DIV[1] _104_ _108_ VGND VGND VPWR VPWR _109_ SKY130_FD_SC_HD__A21OI_2
X_212_ \PLL_CONTRO \PLL_CONTRO _072_ _073_ VGND VGND VPWR VPWR _110_ SKY130_FD_SC_HD__A22O_2
X_213_ \PLL_CONTRO \PLL_CONTRO _088_ _095_ VGND VGND VPWR VPWR _111_ SKY130_FD_SC_HD__O2BB2A_2
X_214_ _110_ _111_ VGND VGND VPWR VPWR _112_ SKY130_FD_SC_HD__OR2_2
X_215_ _110_ _111_ _112_ VGND VGND VPWR VPWR _113_ SKY130_FD_SC_HD__A21BO_2
X_216_ DIV[4] _113_ VGND VGND VPWR VPWR _114_ SKY130_FD_SC_HD__NAND2_2
X_217_ _099_ _101_ _103_ _109_ _114_ VGND VGND VPWR VPWR _115_ SKY130_FD_SC_HD__O221A_2
X_218_ _072_ _073_ DIV[4] _113_ _112_ VGND VGND VPWR VPWR _116_ SKY130_FD_SC_HD__O221AI_2
X_219_ _115_ _116_ VGND VGND VPWR VPWR _117_ SKY130_FD_SC_HD__OR2_2
X_220_ _117_ VGND VGND VPWR VPWR _118_ SKY130_FD_SC_HD__INV_2
X_221_ _081_ _082_ VGND VGND VPWR VPWR _119_ SKY130_FD_SC_HD__OR2_2
X_222_ _119_ VGND VGND VPWR VPWR _120_ SKY130_FD_SC_HD__INV_2
X_223_ _079_ _080_ _119_ VGND VGND VPWR VPWR _015_ SKY130_FD_SC_HD__OR3_2
X_224_ _083_ _084_ _015_ VGND VGND VPWR VPWR _121_ SKY130_FD_SC_HD__OR3_2
X_225_ _085_ _106_ _108_ _102_ _114_ VGND VGND VPWR VPWR _122_ SKY130_FD_SC_HD__O2111AI_2
X_226_ \PLL_CONTRO _087_ \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _123_ SKY130_FD_SC_HD__AND4_2
X_227_ \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _124_ SKY130_FD_SC_HD__OR2_2
X_228_ _124_ VGND VGND VPWR VPWR _125_ SKY130_FD_SC_HD__INV_2
X_229_ \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _126_ SKY130_FD_SC_HD__OR2_2
X_230_ _126_ VGND VGND VPWR VPWR _127_ SKY130_FD_SC_HD__INV_2
X_231_ _124_ _126_ VGND VGND VPWR VPWR _000_ SKY130_FD_SC_HD__OR2_2
X_232_ \PLL_CONTRO _000_ VGND VGND VPWR VPWR _001_ SKY130_FD_SC_HD__OR2_2
X_233_ \PLL_CONTRO \PLL_CONTRO _001_ VGND VGND VPWR VPWR _128_ SKY130_FD_SC_HD__OR3_2
X_234_ _116_ _122_ _117_ _128_ _123_ VGND VGND VPWR VPWR _129_ SKY130_FD_SC_HD__O221A_2
X_235_ _078_ _118_ _121_ _129_ VGND VGND VPWR VPWR _130_ SKY130_FD_SC_HD__O31A_2
X_236_ _130_ VGND VGND VPWR VPWR _131_ SKY130_FD_SC_HD__INV_2
X_237_ \PLL_CONTRO _118_ _083_ _117_ VGND VGND VPWR VPWR _132_ SKY130_FD_SC_HD__A22O_2
X_238_ _083_ _117_ _084_ _132_ VGND VGND VPWR VPWR _133_ SKY130_FD_SC_HD__O22A_2
X_239_ _120_ _125_ VGND VGND VPWR VPWR _134_ SKY130_FD_SC_HD__NOR2_2
X_240_ \PLL_CONTRO _118_ _082_ _117_ VGND VGND VPWR VPWR _135_ SKY130_FD_SC_HD__A22O_2
X_241_ _134_ _135_ _133_ _117_ _125_ VGND VGND VPWR VPWR _136_ SKY130_FD_SC_HD__O32A_2
X_242_ \PLL_CONTRO _118_ _080_ _117_ VGND VGND VPWR VPWR _137_ SKY130_FD_SC_HD__A22O_2
X_243_ _079_ _118_ \PLL_CONTRO _117_ VGND VGND VPWR VPWR _138_ SKY130_FD_SC_HD__O22A_2
X_244_ _138_ VGND VGND VPWR VPWR _139_ SKY130_FD_SC_HD__INV_2
X_245_ _137_ _138_ _136_ _117_ _127_ VGND VGND VPWR VPWR _140_ SKY130_FD_SC_HD__O32A_2
X_246_ _140_ VGND VGND VPWR VPWR _141_ SKY130_FD_SC_HD__INV_2
X_247_ \PLL_CONTRO _118_ _078_ _117_ VGND VGND VPWR VPWR _142_ SKY130_FD_SC_HD__O22A_2
X_248_ _142_ VGND VGND VPWR VPWR _143_ SKY130_FD_SC_HD__INV_2
X_249_ _141_ _142_ _140_ _143_ _131_ VGND VGND VPWR VPWR _144_ SKY130_FD_SC_HD__A221O_2
X_250_ _078_ _130_ _144_ VGND VGND VPWR VPWR _063_ SKY130_FD_SC_HD__O21AI_2
X_251_ _136_ _137_ VGND VGND VPWR VPWR _145_ SKY130_FD_SC_HD__OR2_2
X_252_ _080_ _117_ _145_ VGND VGND VPWR VPWR _146_ SKY130_FD_SC_HD__O21AI_2
X_253_ _146_ VGND VGND VPWR VPWR _147_ SKY130_FD_SC_HD__INV_2
X_254_ _139_ _146_ _138_ _147_ _131_ VGND VGND VPWR VPWR _148_ SKY130_FD_SC_HD__A221O_2
X_255_ _079_ _130_ _148_ VGND VGND VPWR VPWR _062_ SKY130_FD_SC_HD__O21AI_2
X_256_ _136_ _137_ VGND VGND VPWR VPWR _149_ SKY130_FD_SC_HD__NAND2_2
X_257_ _130_ _145_ _149_ \PLL_CONTRO _131_ VGND VGND VPWR VPWR _061_ SKY130_FD_SC_HD__A32O_2
X_258_ _133_ _135_ VGND VGND VPWR VPWR _150_ SKY130_FD_SC_HD__OR2_2
X_259_ \PLL_CONTRO _118_ _133_ VGND VGND VPWR VPWR _151_ SKY130_FD_SC_HD__MUX2_1
X_260_ _082_ _117_ _130_ _151_ VGND VGND VPWR VPWR _152_ SKY130_FD_SC_HD__O211A_2
X_261_ \PLL_CONTRO _152_ \PLL_CONTRO _152_ VGND VGND VPWR VPWR _060_ SKY130_FD_SC_HD__O2BB2A_2
X_262_ _133_ _135_ VGND VGND VPWR VPWR _153_ SKY130_FD_SC_HD__NAND2_2
X_263_ _130_ _150_ _153_ \PLL_CONTRO _131_ VGND VGND VPWR VPWR _059_ SKY130_FD_SC_HD__A32O_2
X_264_ _084_ _132_ _084_ _132_ VGND VGND VPWR VPWR _154_ SKY130_FD_SC_HD__A2BB2O_2
X_265_ _083_ _130_ _131_ _154_ VGND VGND VPWR VPWR _058_ SKY130_FD_SC_HD__O22AI_2
X_266_ \PLL_CONTRO _130_ _084_ _131_ VGND VGND VPWR VPWR _057_ SKY130_FD_SC_HD__O22A_2
X_267_ _075_ _076_ _074_ VGND VGND VPWR VPWR _155_ SKY130_FD_SC_HD__OR3_2
X_268_ _155_ VGND VGND VPWR VPWR _156_ SKY130_FD_SC_HD__INV_2
X_269_ \PLL_CONTRO _156_ VGND VGND VPWR VPWR _157_ SKY130_FD_SC_HD__NAND2_2
X_270_ _072_ _157_ _087_ VGND VGND VPWR VPWR _056_ SKY130_FD_SC_HD__A21OI_2
X_271_ \PLL_CONTRO _156_ \PLL_CONTRO _157_ _086_ VGND VGND VPWR VPWR _055_ SKY130_FD_SC_HD__O221A_2
X_272_ \PLL_CONTRO _156_ \PLL_CONTRO _086_ VGND VGND VPWR VPWR _158_ SKY130_FD_SC_HD__AND4_2
X_273_ _075_ _076_ _074_ VGND VGND VPWR VPWR _159_ SKY130_FD_SC_HD__O21AI_2
X_274_ _086_ _155_ _159_ _158_ VGND VGND VPWR VPWR _054_ SKY130_FD_SC_HD__A31O_2
X_275_ _075_ _076_ \PLL_CONTRO \PLL_CONTRO _086_ VGND VGND VPWR VPWR _160_ SKY130_FD_SC_HD__O221A_2
X_276_ _158_ _160_ VGND VGND VPWR VPWR _053_ SKY130_FD_SC_HD__OR2_2
X_277_ \PLL_CONTRO _156_ \PLL_CONTRO _076_ _087_ VGND VGND VPWR VPWR _052_ SKY130_FD_SC_HD__A311O_2
X_278_ \PLL_CONTRO _126_ VGND VGND VPWR VPWR _004_ SKY130_FD_SC_HD__OR2_2
X_279_ \PLL_CONTRO _004_ VGND VGND VPWR VPWR _007_ SKY130_FD_SC_HD__OR2_2
X_280_ \PLL_CONTRO _080_ VGND VGND VPWR VPWR _161_ SKY130_FD_SC_HD__OR2_2
X_281_ _124_ _161_ \PLL_CONTRO _004_ VGND VGND VPWR VPWR _009_ SKY130_FD_SC_HD__O31A_2
X_282_ \PLL_CONTRO _161_ \PLL_CONTRO _004_ VGND VGND VPWR VPWR _013_ SKY130_FD_SC_HD__O31A_2
X_283_ \PLL_CONTRO _161_ _120_ _004_ VGND VGND VPWR VPWR _006_ SKY130_FD_SC_HD__O31A_2
X_284_ \PLL_CONTRO _161_ _004_ VGND VGND VPWR VPWR _003_ SKY130_FD_SC_HD__O21A_2
X_285_ _079_ \PLL_CONTRO \PLL_CONTRO _124_ _003_ VGND VGND VPWR VPWR _010_ SKY130_FD_SC_HD__O41A_2
X_286_ _079_ \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO _003_ VGND VGND VPWR VPWR _005_ SKY130_FD_SC_HD__O41A_2
X_287_ _079_ \PLL_CONTRO \PLL_CONTRO _120_ _003_ VGND VGND VPWR VPWR _012_ SKY130_FD_SC_HD__O41A_2
X_288_ _120_ _004_ VGND VGND VPWR VPWR _011_ SKY130_FD_SC_HD__OR2_2
X_289_ _079_ \PLL_CONTRO \PLL_CONTRO _003_ VGND VGND VPWR VPWR _002_ SKY130_FD_SC_HD__O31A_2
X_290_ \PLL_CONTRO \PLL_CONTRO _124_ \PLL_CONTRO VGND VGND VPWR VPWR _008_ SKY130_FD_SC_HD__A31O_2
X_291_ \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO \PLL_CONTRO VGND VGND VPWR VPWR _014_ SKY130_FD_SC_HD__A31O_2
X_292_ _078_ _015_ VGND VGND VPWR VPWR _022_ SKY130_FD_SC_HD__NAND2_2
X_293_ \PLL_CONTRO _082_ _126_ \PLL_CONTRO _000_ VGND VGND VPWR VPWR _024_ SKY130_FD_SC_HD__O311A_2
X_294_ _124_ _161_ _078_ VGND VGND VPWR VPWR _162_ SKY130_FD_SC_HD__OR3_2
X_295_ _078_ _126_ _081_ _162_ _024_ VGND VGND VPWR VPWR _017_ SKY130_FD_SC_HD__O311A_2
X_296_ \PLL_CONTRO _082_ _161_ _078_ _017_ VGND VGND VPWR VPWR _025_ SKY130_FD_SC_HD__O41A_2
X_297_ _079_ \PLL_CONTRO _124_ _078_ VGND VGND VPWR VPWR _163_ SKY130_FD_SC_HD__OR4_2
X_298_ _078_ _161_ _081_ _163_ _025_ VGND VGND VPWR VPWR _016_ SKY130_FD_SC_HD__O311A_2
X_299_ _018_ _022_ VGND VGND VPWR VPWR _019_ SKY130_FD_SC_HD__AND2_2
X_300_ _081_ \PLL_CONTRO _078_ _161_ _025_ VGND VGND VPWR VPWR _020_ SKY130_FD_SC_HD__O41A_2
X_301_ _078_ _127_ VGND VGND VPWR VPWR _021_ SKY130_FD_SC_HD__NOR2_2
X_302_ \PLL_CONTRO _126_ _161_ VGND VGND VPWR VPWR _027_ SKY130_FD_SC_HD__AND3_2
X_303_ _079_ \PLL_CONTRO \PLL_CONTRO _027_ VGND VGND VPWR VPWR _023_ SKY130_FD_SC_HD__O31A_2
X_304_ _120_ _125_ _126_ \PLL_CONTRO _000_ VGND VGND VPWR VPWR _028_ SKY130_FD_SC_HD__O311A_2
X_305_ _050_ VGND VGND VPWR VPWR _049_ SKY130_FD_SC_HD__BUF_1
X_306_ _050_ VGND VGND VPWR VPWR _048_ SKY130_FD_SC_HD__BUF_1
X_307_ _050_ VGND VGND VPWR VPWR _047_ SKY130_FD_SC_HD__BUF_1
X_308_ _050_ VGND VGND VPWR VPWR _046_ SKY130_FD_SC_HD__BUF_1
X_309_ _050_ VGND VGND VPWR VPWR _045_ SKY130_FD_SC_HD__BUF_1
X_310_ _050_ VGND VGND VPWR VPWR _044_ SKY130_FD_SC_HD__BUF_1
X_311_ _050_ VGND VGND VPWR VPWR _043_ SKY130_FD_SC_HD__BUF_1
X_312_ _050_ VGND VGND VPWR VPWR _042_ SKY130_FD_SC_HD__BUF_1
X_313_ _050_ VGND VGND VPWR VPWR _041_ SKY130_FD_SC_HD__BUF_1
X_314_ _050_ VGND VGND VPWR VPWR _040_ SKY130_FD_SC_HD__BUF_1
X_315_ _050_ VGND VGND VPWR VPWR _039_ SKY130_FD_SC_HD__BUF_1
X_316_ _050_ VGND VGND VPWR VPWR _038_ SKY130_FD_SC_HD__BUF_1
X_317_ _050_ VGND VGND VPWR VPWR _037_ SKY130_FD_SC_HD__BUF_1
X_318_ _050_ VGND VGND VPWR VPWR _036_ SKY130_FD_SC_HD__BUF_1
X_319_ _050_ VGND VGND VPWR VPWR _035_ SKY130_FD_SC_HD__BUF_1
X_320_ _050_ VGND VGND VPWR VPWR _034_ SKY130_FD_SC_HD__BUF_1
X_321_ _050_ VGND VGND VPWR VPWR _033_ SKY130_FD_SC_HD__BUF_1
X_322_ _050_ VGND VGND VPWR VPWR _032_ SKY130_FD_SC_HD__BUF_1
X_323_ _050_ VGND VGND VPWR VPWR _031_ SKY130_FD_SC_HD__BUF_1
X_324_ _050_ VGND VGND VPWR VPWR _030_ SKY130_FD_SC_HD__BUF_1
X_325_ _050_ VGND VGND VPWR VPWR _029_ SKY130_FD_SC_HD__BUF_1
X_326_ \PLL_CONTRO VGND VGND VPWR VPWR _026_ SKY130_FD_SC_HD__BUF_1
X_327_ _050_ VGND VGND VPWR VPWR _051_ SKY130_FD_SC_HD__BUF_1
X_328_ \PLL_CONTRO VGND VGND VPWR VPWR CLOCKP[0] SKY130_FD_SC_HD__BUF_2
X_329_ _015_ _000_ \PLL_CONTRO VGND VGND VPWR VPWR _018_ SKY130_FD_SC_HD__MUX2_1
X_330_ _012_ EXT_TRIM[11] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_331_ _027_ EXT_TRIM[24] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_332_ _011_ EXT_TRIM[10] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_333_ _026_ EXT_TRIM[23] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_334_ _010_ EXT_TRIM[9] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_335_ _025_ EXT_TRIM[22] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_336_ _009_ EXT_TRIM[8] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_337_ _024_ EXT_TRIM[21] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_338_ _008_ EXT_TRIM[7] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_339_ _023_ EXT_TRIM[20] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_340_ _007_ EXT_TRIM[6] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_341_ _022_ EXT_TRIM[19] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_342_ _006_ EXT_TRIM[5] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_343_ _021_ EXT_TRIM[18] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_344_ _005_ EXT_TRIM[4] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_345_ _020_ EXT_TRIM[17] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_346_ _004_ EXT_TRIM[3] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_347_ _019_ EXT_TRIM[16] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_348_ _003_ EXT_TRIM[2] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_349_ _017_ EXT_TRIM[15] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_350_ _002_ EXT_TRIM[1] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_351_ _016_ EXT_TRIM[14] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_352_ _001_ EXT_TRIM[0] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_353_ _014_ EXT_TRIM[13] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_354_ _013_ EXT_TRIM[12] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_355_ _028_ EXT_TRIM[25] DCO VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__MUX2_1
X_356_ \PLL_CONTRO OSC _029_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_357_ \PLL_CONTRO \PLL_CONTRO _030_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_358_ \PLL_CONTRO \PLL_CONTRO _031_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_359_ \PLL_CONTRO _052_ _032_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_360_ \PLL_CONTRO _053_ _033_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_361_ \PLL_CONTRO _054_ _034_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_362_ \PLL_CONTRO _055_ _035_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_363_ \PLL_CONTRO _056_ _036_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_364_ \PLL_CONTRO _057_ _037_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_365_ \PLL_CONTRO _058_ _038_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_366_ \PLL_CONTRO _059_ _039_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_367_ \PLL_CONTRO _060_ _040_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_368_ \PLL_CONTRO _061_ _041_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_369_ \PLL_CONTRO _062_ _042_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_370_ \PLL_CONTRO _063_ _043_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_371_ \PLL_CONTRO _064_ _044_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_372_ \PLL_CONTRO _065_ _045_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_373_ \PLL_CONTRO _066_ _046_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_374_ \PLL_CONTRO _067_ _047_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_375_ \PLL_CONTRO _068_ _048_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_376_ \PLL_CONTRO _069_ _049_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_377_ \PLL_CONTRO _070_ _050_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X_378_ \PLL_CONTRO _071_ _051_ VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__DFRTP_2
X\RINGOSC.DSTAGE[0].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[0].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[0].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[0].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[0].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[0].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[0].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[10].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[10].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[10].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[10].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[10].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[10].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[10].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[11].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[11].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[11].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[11].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[11].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[11].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[11].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[1].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[1].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[1].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[1].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[1].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[1].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[1].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[2].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[2].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[2].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[2].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[2].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[2].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[2].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[3].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[3].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[3].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[3].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[3].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[3].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[3].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[4].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[4].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[4].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[4].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[4].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[4].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[4].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[5].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[5].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[5].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[5].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[5].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[5].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[5].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[6].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[6].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[6].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[6].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[6].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[6].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[6].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[7].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[7].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[7].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[7].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[7].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[7].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[7].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[8].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[8].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[8].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[8].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[8].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[8].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[8].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.DSTAGE[9].ID.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_2
X\RINGOSC.DSTAGE[9].ID.DELAYBUF1 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.DSTAGE[9].ID.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[9].ID.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.DSTAGE[9].ID.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.DSTAGE[9].ID.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.DSTAGE[9].ID.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.IBUFP00 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_2
X\RINGOSC.IBUFP01 \RINGOS VGND VGND VPWR VPWR \PLL_CONTRO SKY130_FD_SC_HD__CLKINV_8
X\RINGOSC.IBUFP10 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_2
X\RINGOSC.IBUFP11 \RINGOS VGND VGND VPWR VPWR CLOCKP[1] SKY130_FD_SC_HD__CLKINV_8
X\RINGOSC.ISS.CONST1 VPB VNB VPWR VGND \RINGOS SKY130_FD_SC_HD__CONB_1
X\RINGOSC.ISS.CTRLEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__OR2_2
X\RINGOSC.ISS.DELAYBUF0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKBUF_1
X\RINGOSC.ISS.DELAYEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.ISS.DELAYEN1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_2
X\RINGOSC.ISS.DELAYENB0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_8
X\RINGOSC.ISS.DELAYENB1 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVN_4
X\RINGOSC.ISS.DELAYINT0 \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__CLKINV_1
X\RINGOSC.ISS.RESETEN0 \RINGOS \RINGOS VGND VGND VPWR VPWR \RINGOS SKY130_FD_SC_HD__EINVP_1

.ENDS DIGITAL_PLL