* Extracted by KLayout on : 22/12/2021 04:25

.SUBCKT digital_pll osc clockp[0] clockp[1] div[0] VPWR div[1] div[2]
+ ext_trim[24] div[3] div[4] ext_trim[23] resetb enable dco ext_trim[0]
+ ext_trim[25] ext_trim[1] ext_trim[13] ext_trim[22] ext_trim[11] ext_trim[12]
+ ext_trim[14] ext_trim[2] ext_trim[21] ext_trim[18] ext_trim[10] ext_trim[9]
+ ext_trim[3] ext_trim[15] ext_trim[5] ext_trim[19] ext_trim[20] ext_trim[4]
+ ext_trim[6] ext_trim[17] ext_trim[16] ext_trim[7] ext_trim[8] VGND
X$1 VPWR osc VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$2 VGND \$25 \$14 \$12 osc VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$3 VPWR VGND clockp[0] VPWR \$12 VGND sky130_fd_sc_hd__buf_2
X$4 VPWR VGND \$11 VPWR \$4 \$9 VGND sky130_fd_sc_hd__nor2_2
X$5 VPWR VPWR \$11 \$29 \$9 VGND \$4 VGND sky130_fd_sc_hd__a21oi_2
X$6 VGND \$96 \$9 \$11 \$49 \$4 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$7 VPWR \$18 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$8 VGND \$5 \$71 \$12 \$73 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$9 VPWR VGND dco VPWR \$5 \$164 VGND sky130_fd_sc_hd__nor2_2
X$10 VPWR \$52 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$11 VPWR \$94 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$12 VPWR \$50 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$13 VPWR \$95 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$14 VPWR \$7 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$15 VPWR \$121 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$16 VPWR \$143 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$17 VPWR \$142 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$18 VPWR \$67 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$19 VPWR \$133 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$20 VPWR \$132 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$21 VPWR \$32 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$22 VPWR \$25 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$23 VPWR \$35 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$24 VPWR \$65 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$25 VPWR \$80 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$26 VPWR \$147 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$27 VPWR \$24 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$28 VPWR \$150 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$29 VPWR \$23 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$30 VPWR \$106 VGND VPWR \$5 VGND sky130_fd_sc_hd__buf_1
X$31 VGND clockp[1] \$169 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$32 VGND \$7 \$11 \$12 \$53 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$33 VGND \$37 \$63 \$64 \$31 \$8 VPWR VPWR VGND sky130_fd_sc_hd__and4_2
X$34 VGND \$24 \$8 \$12 \$16 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$35 VPWR \$16 VPWR VGND \$37 \$8 VGND sky130_fd_sc_hd__or2_2
X$36 VGND \$8 \$31 \$30 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$37 VGND \$11 \$9 \$19 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$38 VGND \$18 \$9 \$12 \$19 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$39 VPWR \$36 VPWR VGND \$20 \$10 \$21 VGND sky130_fd_sc_hd__or3_2
X$40 VPWR VGND VPWR \$10 \$15 VGND sky130_fd_sc_hd__inv_2
X$41 VGND \$27 \$15 \$45 \$21 \$10 \$13 VPWR VPWR VGND sky130_fd_sc_hd__o221a_2
X$42 VPWR \$10 VGND \$21 \$60 VPWR \$36 VGND sky130_fd_sc_hd__o21ai_2
X$43 VPWR VGND VPWR \$36 \$11 VGND sky130_fd_sc_hd__inv_2
X$44 VGND \$35 \$38 \$12 \$14 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$45 VGND \$12 \$139 VPWR VPWR VGND sky130_fd_sc_hd__clkinv_8
X$46 VGND \$147 \$113 \$12 \$108 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$47 VGND \$143 \$144 \$12 \$137 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$48 VGND \$94 \$45 \$12 \$89 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$49 VGND \$23 \$15 \$12 \$22 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$50 VGND \$95 \$82 \$12 \$81 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$51 VGND \$80 \$77 \$12 \$104 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$52 VGND \$150 \$158 \$12 \$146 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$53 VGND \$65 \$42 \$12 \$38 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$54 VGND \$106 \$70 \$12 \$110 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$55 VGND \$50 \$34 \$12 \$51 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$56 VGND \$67 \$75 \$12 \$74 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$57 VGND \$142 \$166 \$12 \$165 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$58 VGND \$32 \$31 \$12 \$30 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$59 VGND \$52 \$63 \$12 \$56 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$60 VGND \$133 \$131 \$12 \$130 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$61 VGND \$121 \$126 \$12 \$115 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$62 VGND \$132 \$97 \$12 \$120 VPWR VPWR VGND sky130_fd_sc_hd__dfrtp_2
X$63 VPWR \$22 VPWR VGND \$13 \$62 VGND sky130_fd_sc_hd__or2_2
X$64 VGND \$41 \$34 \$15 \$34 \$15 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$65 VGND \$15 \$34 \$51 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$66 VGND \$46 \$15 \$44 \$41 \$34 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$67 VGND \$39 div[0] \$43 \$33 div[1] \$47 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$68 VPWR VGND VPWR \$59 div[0] VGND sky130_fd_sc_hd__inv_2
X$69 VPWR div[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$70 VPWR div[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$71 VPWR \$53 VPWR VGND \$60 \$20 \$27 \$62 VGND sky130_fd_sc_hd__a31o_2
X$72 VPWR VGND VPWR \$55 \$20 VGND sky130_fd_sc_hd__inv_2
X$73 VGND \$89 \$97 \$55 \$70 \$21 \$37 VPWR VPWR VGND sky130_fd_sc_hd__a311o_2
X$74 VPWR VPWR \$21 \$40 \$61 VGND \$46 VGND sky130_fd_sc_hd__a21oi_2
X$75 VPWR VGND VPWR \$21 \$45 VGND sky130_fd_sc_hd__inv_2
X$76 VPWR VGND \$21 VPWR \$46 \$61 VGND sky130_fd_sc_hd__nor2_2
X$77 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$78 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$79 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$80 VPWR \$312 VPWR \$283 VGND \$317 VGND sky130_fd_sc_hd__einvp_2
X$81 VPWR \$288 VPWR \$287 VGND \$315 VGND sky130_fd_sc_hd__einvp_2
X$82 VPWR \$315 VGND VPWR \$289 VGND sky130_fd_sc_hd__clkbuf_1
X$83 VPWR VPWR VGND \$317 \$288 VGND sky130_fd_sc_hd__clkinv_1
X$84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$85 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$86 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$87 VPWR \$295 VPWR \$301 VGND \$318 VGND sky130_fd_sc_hd__einvp_2
X$88 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$89 VPWR \$316 VPWR \$310 VGND \$313 VGND sky130_fd_sc_hd__einvp_2
X$90 VPWR VPWR VGND \$318 \$316 VGND sky130_fd_sc_hd__clkinv_1
X$91 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$93 VPWR ext_trim[8] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$94 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$95 VPWR ext_trim[7] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$96 VGND \$311 ext_trim[7] \$220 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$97 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$99 VPWR \$314 VPWR \$311 VGND \$282 VGND sky130_fd_sc_hd__einvp_2
X$100 VPWR \$286 VPWR \$302 VGND \$303 VGND sky130_fd_sc_hd__einvp_2
X$101 VGND \$310 ext_trim[17] \$240 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$102 VPWR ext_trim[17] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$103 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$105 VGND \$287 ext_trim[16] \$276 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$106 VPWR \$309 VPWR \$306 VGND \$305 VGND sky130_fd_sc_hd__einvp_2
X$107 VPWR ext_trim[16] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$108 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$109 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$110 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$111 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$112 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$113 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$114 VPWR VGND VPWR \$43 \$40 VGND sky130_fd_sc_hd__inv_2
X$115 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$116 VGND \$48 \$44 \$29 \$44 VPWR \$29 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$118 VGND \$46 \$41 \$33 \$46 \$41 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2ai_2
X$119 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$121 VPWR VGND VPWR \$37 \$27 VGND sky130_fd_sc_hd__inv_2
X$122 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$123 VGND \$27 \$38 \$42 \$38 VPWR \$42 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$124 VPWR \$I1325 VGND VPWR sky130_fd_sc_hd__fill_2
X$125 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$126 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$127 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$128 VPWR VPWR \$39 \$33 VGND div[1] VGND sky130_fd_sc_hd__nand2_2
X$129 VGND \$57 \$54 \$58 \$47 \$40 \$59 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2111ai_2
X$130 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$131 VPWR \$I1346 VGND VPWR sky130_fd_sc_hd__fill_2
X$132 VPWR VGND VPWR \$49 \$44 VGND sky130_fd_sc_hd__inv_2
X$133 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$134 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$135 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$137 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$138 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$139 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$140 VGND \$63 \$31 \$56 \$27 \$37 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$141 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$143 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$144 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$145 VPWR div[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$146 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$147 VPWR \$69 VPWR \$66 VGND \$48 div[2] \$58 VGND sky130_fd_sc_hd__o211a_2
X$148 VPWR VPWR div[1] \$78 \$33 VGND \$47 VGND sky130_fd_sc_hd__a21oi_2
X$149 VGND \$70 \$71 \$73 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$151 VGND \$55 \$97 \$62 \$70 \$27 VPWR VPWR VGND sky130_fd_sc_hd__and4_2
X$152 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$153 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$155 VGND \$81 \$72 \$123 \$76 \$82 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$156 VPWR \$182 VPWR VGND \$79 \$77 \$82 VGND sky130_fd_sc_hd__or3_2
X$157 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$158 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$159 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$160 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$161 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$162 VPWR div[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$163 VPWR div[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$164 VGND \$57 \$84 \$78 \$87 \$69 \$86 VPWR VPWR VGND sky130_fd_sc_hd__o221a_2
X$165 VPWR VGND VPWR \$84 \$58 VGND sky130_fd_sc_hd__inv_2
X$166 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$167 VPWR VGND \$70 VPWR \$88 \$71 VGND sky130_fd_sc_hd__nor2_2
X$168 VPWR VPWR VGND \$100 \$88 \$70 \$71 VGND sky130_fd_sc_hd__a21o_2
X$169 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$171 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$172 VGND \$45 \$75 \$74 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$173 VPWR VGND VPWR \$61 \$75 VGND sky130_fd_sc_hd__inv_2
X$174 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$175 VGND \$64 \$101 \$79 \$54 \$91 \$92 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$176 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$177 VGND \$93 \$77 \$85 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$179 VPWR \$I1345 VGND VPWR sky130_fd_sc_hd__fill_2
X$180 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$181 VPWR ext_trim[2] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$182 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$183 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$184 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$185 VPWR VPWR VGND \$216 \$238 VGND sky130_fd_sc_hd__clkbuf_2
X$186 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$187 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$189 VPWR VPWR VGND \$213 \$218 VGND sky130_fd_sc_hd__clkinv_1
X$190 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$191 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$192 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$193 VGND \$184 ext_trim[12] \$234 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$194 VGND \$290 \$214 \$158 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$195 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$196 VGND \$239 \$214 \$205 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$197 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$198 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$199 VGND \$219 ext_trim[14] \$235 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$201 VGND \$235 \$111 \$221 \$236 \$230 \$233 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$202 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$203 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$204 VGND \$240 \$233 \$221 \$111 \$131 \$236 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$205 VPWR \$111 VPWR VGND \$241 \$205 \$221 VGND sky130_fd_sc_hd__or3_2
X$206 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$207 VPWR ext_trim[21] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$208 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$209 VPWR VPWR VGND \$232 \$207 VGND sky130_fd_sc_hd__clkbuf_2
X$210 VGND \$243 ext_trim[22] \$233 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$211 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$212 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$213 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$214 VGND \$258 ext_trim[2] \$214 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$215 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$216 VGND \$238 \$248 \$245 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$217 VPWR \$259 VGND VPWR \$238 VGND sky130_fd_sc_hd__clkbuf_1
X$218 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$219 VPWR VPWR VGND \$260 \$249 VGND sky130_fd_sc_hd__clkinv_1
X$220 VGND \$246 \$249 \$247 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$221 VGND \$234 \$126 \$221 \$158 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$223 VPWR \$250 VPWR VGND \$244 \$158 VGND sky130_fd_sc_hd__or2_2
X$224 VGND \$261 \$205 \$221 \$126 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$225 VGND \$226 ext_trim[10] \$251 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$226 VPWR \$251 VPWR VGND \$244 \$190 VGND sky130_fd_sc_hd__or2_2
X$227 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$228 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$229 VPWR ext_trim[14] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$230 VGND \$233 \$252 \$111 \$221 \$153 \$158 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$231 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$232 VGND \$254 \$158 \$153 \$187 \$126 \$204 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$233 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$235 VGND \$262 ext_trim[21] \$254 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$236 VPWR \$232 VPWR \$271 VGND \$255 VGND sky130_fd_sc_hd__einvp_2
X$237 VPWR \$256 VPWR \$243 VGND \$257 VGND sky130_fd_sc_hd__einvp_2
X$238 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$239 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$240 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$241 VGND \$289 \$283 \$312 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$242 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$243 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$244 VGND \$289 \$288 \$287 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$245 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$246 VPWR VPWR VGND \$312 \$307 VGND sky130_fd_sc_hd__clkbuf_2
X$247 VPWR VPWR VGND \$273 \$289 VGND sky130_fd_sc_hd__clkbuf_2
X$248 VGND \$307 \$301 \$295 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$249 VPWR ext_trim[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$251 VGND \$301 ext_trim[4] \$290 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$252 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$253 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$254 VPWR VPWR VGND \$295 \$246 VGND sky130_fd_sc_hd__clkbuf_2
X$255 VGND \$307 \$316 \$310 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$256 VPWR ext_trim[6] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$257 VGND \$299 ext_trim[6] \$250 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$258 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$260 VGND \$269 \$299 \$300 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$261 VPWR \$313 VGND VPWR \$307 VGND sky130_fd_sc_hd__clkbuf_1
X$262 VGND \$306 ext_trim[8] \$261 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$263 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$264 VPWR VPWR VGND \$300 \$308 VGND sky130_fd_sc_hd__clkbuf_2
X$265 VPWR \$300 VPWR \$299 VGND \$291 VGND sky130_fd_sc_hd__einvp_2
X$266 VGND \$308 \$311 \$314 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$267 VPWR VPWR VGND \$291 \$284 VGND sky130_fd_sc_hd__clkinv_1
X$268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$269 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$270 VGND \$302 ext_trim[20] \$229 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$271 VGND \$308 \$286 \$302 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$272 VPWR \$303 VGND VPWR \$308 VGND sky130_fd_sc_hd__clkbuf_1
X$273 VPWR ext_trim[20] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$274 VGND \$281 ext_trim[19] \$267 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$275 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$276 VPWR \$293 VPWR \$262 VGND \$304 VGND sky130_fd_sc_hd__einvp_2
X$277 VPWR ext_trim[19] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$279 VPWR \$I1205 VGND VPWR sky130_fd_sc_hd__fill_1
X$280 VGND \$294 \$293 \$262 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$281 VPWR VPWR VGND \$314 \$294 VGND sky130_fd_sc_hd__clkbuf_2
X$282 VGND \$294 \$306 \$309 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$283 VPWR \$304 VGND VPWR \$294 VGND sky130_fd_sc_hd__clkbuf_1
X$284 VPWR VPWR VGND \$305 \$293 VGND sky130_fd_sc_hd__clkinv_1
X$285 VPWR VPWR VGND \$309 \$268 VGND sky130_fd_sc_hd__clkbuf_2
X$286 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$287 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$288 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$289 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$290 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$291 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$292 VPWR ext_trim[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$293 VGND \$197 ext_trim[0] \$182 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$294 VGND \$202 \$197 \$183 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$295 VPWR \$183 VPWR \$197 VGND \$175 VGND sky130_fd_sc_hd__einvp_2
X$296 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$297 VPWR \$176 VPWR \$193 VGND \$192 VGND sky130_fd_sc_hd__einvp_2
X$298 VGND \$202 \$176 \$193 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$299 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$301 VPWR VPWR \$181 VGND \$164 \$198 VGND sky130_fd_sc_hd__einvp_1
X$302 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$303 VPWR \$199 VPWR VGND \$184 \$164 VGND sky130_fd_sc_hd__or2_2
X$304 VGND \$171 \$199 \$181 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$305 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$306 VPWR \$181 VPWR \$184 VGND \$194 VGND sky130_fd_sc_hd__einvp_2
X$307 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$308 VGND \$171 \$185 \$186 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$309 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$311 VPWR VPWR VGND \$194 \$185 VGND sky130_fd_sc_hd__clkinv_1
X$312 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$313 VPWR \$185 VPWR \$186 VGND \$177 VGND sky130_fd_sc_hd__einvp_2
X$314 VGND \$193 ext_trim[13] \$203 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$315 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$316 VPWR \$195 VGND \$101 \$155 VPWR \$178 VGND sky130_fd_sc_hd__o21ai_2
X$317 VPWR \$203 VPWR VGND \$158 \$166 \$144 \$126 VGND sky130_fd_sc_hd__a31o_2
X$318 VPWR VGND VPWR \$156 \$144 VGND sky130_fd_sc_hd__inv_2
X$319 VPWR \$187 VPWR VGND \$166 \$144 VGND sky130_fd_sc_hd__or2_2
X$320 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$321 VPWR VGND VPWR \$161 \$187 VGND sky130_fd_sc_hd__inv_2
X$322 VPWR VGND VPWR \$195 \$166 VGND sky130_fd_sc_hd__inv_2
X$323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$324 VGND \$186 ext_trim[25] \$188 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$325 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$326 VGND \$188 \$190 \$172 \$187 \$126 \$204 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$327 VPWR VGND \$190 VPWR \$170 \$172 VGND sky130_fd_sc_hd__nor2_2
X$328 VPWR \$182 VPWR VGND \$204 \$126 VGND sky130_fd_sc_hd__or2_2
X$329 VPWR ext_trim[25] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$330 VPWR \$I1211 VGND VPWR sky130_fd_sc_hd__fill_1
X$331 VPWR VGND VPWR \$111 \$126 VGND sky130_fd_sc_hd__inv_2
X$332 VPWR VGND VPWR \$172 \$205 VGND sky130_fd_sc_hd__inv_2
X$333 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$334 VPWR \$171 VPWR \$206 VGND \$200 VGND sky130_fd_sc_hd__einvp_2
X$335 VPWR VPWR VGND \$200 \$191 VGND sky130_fd_sc_hd__clkinv_1
X$336 VPWR \$191 VPWR \$180 VGND \$179 VGND sky130_fd_sc_hd__einvp_2
X$337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$338 VGND \$174 \$206 \$171 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$339 VGND \$174 \$191 \$180 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$340 VPWR \$201 VPWR \$168 VGND \$196 VGND sky130_fd_sc_hd__einvp_2
X$341 VPWR \$196 VGND VPWR \$207 VGND sky130_fd_sc_hd__clkbuf_1
X$342 VPWR ext_trim[23] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$343 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$344 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$345 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$346 VPWR \$I1207 VGND VPWR sky130_fd_sc_hd__fill_1
X$347 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$348 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$349 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$351 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$352 VPWR \$I1214 VGND VPWR sky130_fd_sc_hd__fill_1
X$353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$354 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$355 VPWR \$I1212 VGND VPWR sky130_fd_sc_hd__fill_1
X$356 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$357 VPWR \$I1324 VGND VPWR sky130_fd_sc_hd__fill_2
X$358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$359 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$360 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$362 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$363 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$364 VPWR div[1] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$365 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$367 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$368 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$370 VPWR \$I1325 VGND VPWR sky130_fd_sc_hd__fill_2
X$371 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$372 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$373 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$374 VGND \$283 ext_trim[3] \$244 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$375 VPWR ext_trim[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$376 VGND \$238 \$258 \$273 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$377 VPWR \$273 VPWR \$258 VGND \$277 VGND sky130_fd_sc_hd__einvp_2
X$378 VPWR \$248 VPWR \$245 VGND \$259 VGND sky130_fd_sc_hd__einvp_2
X$379 VPWR VPWR VGND \$277 \$248 VGND sky130_fd_sc_hd__clkinv_1
X$380 VPWR ext_trim[5] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$381 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$382 VPWR \$I1259 VGND VPWR sky130_fd_sc_hd__fill_1
X$383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$384 VGND \$265 ext_trim[5] \$278 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$385 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$386 VGND \$246 \$265 \$274 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$387 VPWR \$274 VPWR \$265 VGND \$260 VGND sky130_fd_sc_hd__einvp_2
X$388 VPWR \$249 VPWR \$247 VGND \$279 VGND sky130_fd_sc_hd__einvp_2
X$389 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$390 VGND \$278 \$126 \$221 \$190 \$244 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$391 VPWR \$279 VGND VPWR \$246 VGND sky130_fd_sc_hd__clkbuf_1
X$392 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$394 VPWR VGND VPWR \$214 \$244 \$221 \$126 VGND sky130_fd_sc_hd__o21a_2
X$395 VGND \$271 ext_trim[9] \$239 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$396 VPWR VPWR VGND \$274 \$269 VGND sky130_fd_sc_hd__clkbuf_2
X$397 VPWR ext_trim[10] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$398 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$399 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$400 VGND \$269 \$284 \$281 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$401 VPWR ext_trim[9] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$402 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$403 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$404 VPWR \$275 VGND VPWR \$269 VGND sky130_fd_sc_hd__clkbuf_1
X$405 VPWR VGND \$111 VPWR \$264 \$161 VGND sky130_fd_sc_hd__nor2_2
X$406 VPWR \$284 VPWR \$281 VGND \$275 VGND sky130_fd_sc_hd__einvp_2
X$407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$408 VGND \$247 ext_trim[18] \$264 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$409 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$410 VGND \$245 ext_trim[15] \$252 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$411 VPWR ext_trim[18] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$412 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$413 VPWR VPWR VGND \$282 \$286 VGND sky130_fd_sc_hd__clkinv_1
X$414 VGND \$252 \$111 \$187 \$236 \$241 \$254 VPWR VPWR VGND
+ sky130_fd_sc_hd__o311a_2
X$415 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$416 VGND \$270 \$204 \$117 \$126 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$417 VPWR VPWR \$270 \$267 \$276 VGND VGND sky130_fd_sc_hd__and2_2
X$418 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$419 VPWR \$I1209 VGND VPWR sky130_fd_sc_hd__fill_1
X$420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$421 VPWR VPWR \$267 \$117 VGND \$111 VGND sky130_fd_sc_hd__nand2_2
X$422 VGND \$268 \$271 \$232 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$423 VPWR ext_trim[15] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$424 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$425 VPWR VPWR VGND \$255 \$256 VGND sky130_fd_sc_hd__clkinv_1
X$426 VGND \$268 \$256 \$243 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$427 VPWR \$257 VGND VPWR \$268 VGND sky130_fd_sc_hd__clkbuf_1
X$428 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$429 VPWR \$I1260 VGND VPWR sky130_fd_sc_hd__fill_1
X$430 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$431 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$432 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$433 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$434 VPWR ext_trim[0] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$435 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$436 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$437 VPWR div[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$438 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$439 VPWR \$169 \$274 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$440 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$441 VPWR VPWR VGND \$175 \$176 VGND sky130_fd_sc_hd__clkinv_1
X$442 VPWR VGND VPWR \$114 \$113 VGND sky130_fd_sc_hd__inv_2
X$443 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$444 VPWR resetb VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$445 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$446 VPWR \$I1236 VGND VPWR sky130_fd_sc_hd__fill_1
X$447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$448 VPWR VPWR \$164 resetb VGND enable VGND sky130_fd_sc_hd__nand2_2
X$449 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$450 VPWR enable VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$451 VPWR \$139 \$181 VPWR VGND VGND sky130_fd_sc_hd__clkinv_2
X$452 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$453 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$454 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$456 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$457 VPWR \$177 VGND VPWR \$171 VGND sky130_fd_sc_hd__clkbuf_1
X$458 VPWR VGND VPWR \$160 \$155 VGND sky130_fd_sc_hd__inv_2
X$459 VPWR \$156 VGND \$76 \$137 VPWR \$167 VGND sky130_fd_sc_hd__o21ai_2
X$460 VPWR VGND VPWR \$152 \$151 VGND sky130_fd_sc_hd__inv_2
X$461 VGND \$151 \$152 \$167 \$123 \$160 \$155 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_2
X$462 VGND \$165 \$76 \$178 \$123 \$166 \$134 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$463 VGND \$151 \$144 \$101 \$102 \$156 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$464 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$465 VGND \$195 \$166 \$141 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$467 VGND \$124 \$141 \$151 \$140 \$161 \$101 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$468 VPWR \$178 VPWR VGND \$141 \$140 VGND sky130_fd_sc_hd__or2_2
X$469 VGND \$140 \$170 \$138 \$118 \$172 \$101 VPWR VPWR VGND
+ sky130_fd_sc_hd__o32a_2
X$470 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$471 VGND \$153 \$131 \$138 \$101 \$102 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$472 VPWR \$I1211 VGND VPWR sky130_fd_sc_hd__fill_1
X$473 VGND \$157 \$102 \$131 \$118 VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$474 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$475 VPWR \$157 VPWR \$76 VGND \$101 \$153 \$149 VGND sky130_fd_sc_hd__o211a_2
X$476 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$478 VPWR VGND VPWR \$153 \$131 VGND sky130_fd_sc_hd__inv_2
X$479 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$480 VGND \$146 \$149 \$158 \$149 \$158 VPWR VPWR VGND
+ sky130_fd_sc_hd__o2bb2a_2
X$481 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$482 VPWR \$179 VGND VPWR \$174 VGND sky130_fd_sc_hd__clkbuf_1
X$483 VGND \$180 ext_trim[24] \$173 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$484 VGND \$168 ext_trim[23] \$159 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$485 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$486 VPWR \$159 VGND VPWR \$126 VGND sky130_fd_sc_hd__buf_1
X$487 VPWR ext_trim[24] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$488 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$489 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$490 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$491 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$492 VPWR div[4] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$493 VPWR div[3] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$494 VPWR VPWR \$57 \$119 VGND div[4] VGND sky130_fd_sc_hd__nand2_2
X$495 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$496 VGND \$112 \$91 div[4] \$119 \$122 \$114 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221ai_2
X$497 VPWR \$112 VPWR VGND \$105 \$107 VGND sky130_fd_sc_hd__or2_2
X$498 VPWR \$I1236 VGND VPWR sky130_fd_sc_hd__fill_1
X$499 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$500 VPWR VGND VPWR \$122 \$97 VGND sky130_fd_sc_hd__inv_2
X$501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$502 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$503 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$504 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$505 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$507 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$508 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$509 VPWR VGND VPWR \$123 \$76 VGND sky130_fd_sc_hd__inv_2
X$510 VPWR VGND VPWR \$127 \$124 VGND sky130_fd_sc_hd__inv_2
X$511 VGND \$128 \$111 \$101 \$102 \$126 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$512 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$513 VPWR VGND VPWR \$129 \$128 VGND sky130_fd_sc_hd__inv_2
X$514 VPWR VPWR \$134 \$141 VGND \$140 VGND sky130_fd_sc_hd__nand2_2
X$515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$516 VGND \$124 \$127 \$116 \$123 \$129 \$128 VPWR VPWR VGND
+ sky130_fd_sc_hd__a221o_2
X$517 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$518 VPWR VPWR \$135 \$138 VGND \$118 VGND sky130_fd_sc_hd__nand2_2
X$519 VGND \$130 \$76 \$145 \$123 \$131 \$135 VPWR VPWR VGND
+ sky130_fd_sc_hd__a32o_2
X$520 VPWR \$145 VPWR VGND \$138 \$118 VGND sky130_fd_sc_hd__or2_2
X$521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$522 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$523 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$524 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$525 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$526 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$527 VGND \$48 div[2] \$69 div[3] \$99 VPWR VPWR VGND sky130_fd_sc_hd__a22oi_2
X$528 VPWR VGND VPWR \$87 \$66 VGND sky130_fd_sc_hd__inv_2
X$529 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$530 VGND \$99 \$100 \$96 \$100 VPWR \$96 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$531 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$533 VGND \$105 \$71 \$70 \$96 \$88 VPWR VPWR VGND sky130_fd_sc_hd__o2bb2a_2
X$534 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$535 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$536 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$537 VPWR \$101 VPWR VGND \$91 \$86 VGND sky130_fd_sc_hd__or2_2
X$538 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$539 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$541 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$542 VPWR VGND VPWR \$72 \$82 VGND sky130_fd_sc_hd__inv_2
X$543 VGND \$76 \$111 \$102 \$103 \$92 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$544 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$545 VGND \$123 \$104 \$98 \$76 \$93 VPWR VPWR VGND sky130_fd_sc_hd__o22ai_2
X$546 VGND \$98 \$72 \$85 \$72 VPWR \$85 VPWR VGND sky130_fd_sc_hd__a2bb2o_2
X$547 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$548 VPWR \$I1345 VGND VPWR sky130_fd_sc_hd__fill_2
X$549 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$550 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$551 VPWR \$66 VPWR VGND \$99 div[3] VGND sky130_fd_sc_hd__or2_2
X$552 VPWR VPWR VGND \$119 \$112 \$107 \$105 VGND sky130_fd_sc_hd__a21bo_2
X$553 VGND \$122 \$97 \$107 \$114 \$113 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$554 VGND \$97 \$113 \$108 \$37 \$27 VPWR VPWR VGND sky130_fd_sc_hd__a22o_2
X$555 VPWR VPWR \$122 \$120 \$109 VGND \$37 VGND sky130_fd_sc_hd__a21oi_2
X$556 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$557 VGND \$27 \$97 \$109 \$55 \$70 \$110 VPWR VPWR VGND
+ sky130_fd_sc_hd__o221a_2
X$558 VPWR VPWR \$109 \$55 VGND \$70 VGND sky130_fd_sc_hd__nand2_2
X$559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$560 VPWR VGND VPWR \$102 \$101 VGND sky130_fd_sc_hd__inv_2
X$561 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$562 VPWR \$111 VGND \$76 \$115 VPWR \$116 VGND sky130_fd_sc_hd__o21ai_2
X$563 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_6
X$564 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$565 VPWR \$117 VPWR VGND \$103 \$93 \$72 VGND sky130_fd_sc_hd__or3_2
X$566 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$567 VGND \$118 \$72 \$85 \$101 \$93 VPWR VPWR VGND sky130_fd_sc_hd__o22a_2
X$568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$569 VPWR VGND VPWR \$93 \$77 VGND sky130_fd_sc_hd__inv_2
X$570 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$571 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$572 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$573 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$574 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$575 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$576 VGND \$223 ext_trim[1] \$212 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$577 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$578 VPWR \$216 VPWR \$223 VGND \$213 VGND sky130_fd_sc_hd__einvp_2
X$579 VPWR VPWR VGND \$183 \$224 VGND sky130_fd_sc_hd__clkbuf_2
X$580 VPWR \$192 VGND VPWR \$202 VGND sky130_fd_sc_hd__clkbuf_1
X$581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$582 VPWR \$218 VPWR \$219 VGND \$217 VGND sky130_fd_sc_hd__einvp_2
X$583 VPWR VPWR VGND \$181 \$202 VGND sky130_fd_sc_hd__clkbuf_2
X$584 VPWR VPWR VGND \$198 VGND sky130_fd_sc_hd__conb_1
X$585 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_12
X$586 VGND \$212 \$156 \$166 \$126 \$214 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$587 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$588 VPWR \$220 VPWR VGND \$205 \$166 \$144 \$126 VGND sky130_fd_sc_hd__a31o_2
X$589 VPWR \$221 VPWR VGND \$195 \$144 VGND sky130_fd_sc_hd__or2_2
X$590 VPWR ext_trim[13] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$591 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$593 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$594 VPWR \$211 VPWR VGND \$117 \$156 \$195 VGND sky130_fd_sc_hd__or3_2
X$595 VPWR \$211 VPWR VGND \$153 \$236 VGND sky130_fd_sc_hd__or2_2
X$596 VPWR VGND VPWR \$190 \$211 VGND sky130_fd_sc_hd__inv_2
X$597 VPWR \$126 \$187 \$221 VGND VPWR \$173 VGND sky130_fd_sc_hd__and3_2
X$598 VPWR \$205 VPWR VGND \$131 \$158 VGND sky130_fd_sc_hd__or2_2
X$599 VPWR \$I1336 VGND VPWR sky130_fd_sc_hd__fill_2
X$600 VPWR VPWR VGND \$215 \$174 VGND sky130_fd_sc_hd__clkbuf_2
X$601 VPWR \$215 VPWR \$226 VGND \$222 VGND sky130_fd_sc_hd__einvp_2
X$602 VGND \$207 \$201 \$168 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$603 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$604 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$605 VPWR dco VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$606 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$607 VGND \$224 \$223 \$216 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$608 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$609 VGND \$224 \$218 \$219 VPWR VPWR VGND sky130_fd_sc_hd__einvn_4
X$610 VPWR \$217 VGND VPWR \$224 VGND sky130_fd_sc_hd__clkbuf_1
X$611 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_1
X$612 VGND \$206 ext_trim[11] \$225 dco VPWR VPWR VGND sky130_fd_sc_hd__mux2_1
X$613 VPWR ext_trim[11] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$614 VPWR ext_trim[12] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$615 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$617 VGND \$225 \$214 \$190 \$126 \$166 \$156 VPWR VPWR VGND
+ sky130_fd_sc_hd__o41a_2
X$618 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_4
X$619 VPWR \$244 VPWR VGND \$187 \$126 VGND sky130_fd_sc_hd__or2_2
X$620 VPWR VGND VGND VPWR sky130_fd_sc_hd__fill_2
X$621 VPWR \$205 \$166 VGND \$156 VPWR \$230 \$111 VGND sky130_fd_sc_hd__or4_2
X$622 VGND \$229 \$156 \$166 \$158 \$173 VPWR VPWR VGND sky130_fd_sc_hd__o31a_2
X$623 VPWR VPWR VGND VGND sky130_fd_sc_hd__decap_8
X$624 VPWR \$204 VPWR VGND \$187 \$205 VGND sky130_fd_sc_hd__or2_2
X$625 VPWR VGND VPWR \$236 \$158 VGND sky130_fd_sc_hd__inv_2
X$626 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
X$627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X$628 VGND \$207 \$226 \$215 VPWR VPWR VGND sky130_fd_sc_hd__einvn_8
X$629 VPWR VPWR VGND \$222 \$201 VGND sky130_fd_sc_hd__clkinv_1
X$630 VPWR ext_trim[22] VPWR VGND VGND sky130_fd_sc_hd__diode_2
X$631 VPWR VGND VPWR VGND sky130_fd_sc_hd__decap_3
.ENDS digital_pll

.SUBCKT sky130_fd_sc_hd__o22a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22a_2

.SUBCKT sky130_fd_sc_hd__o22ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o22ai_2

.SUBCKT sky130_fd_sc_hd__and4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__and4_2

.SUBCKT sky130_fd_sc_hd__o2bb2ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o2bb2ai_2

.SUBCKT sky130_fd_sc_hd__o211a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o211a_2

.SUBCKT sky130_fd_sc_hd__o2111ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o2111ai_2

.SUBCKT sky130_fd_sc_hd__buf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_2

.SUBCKT sky130_fd_sc_hd__o221ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221ai_2

.SUBCKT sky130_fd_sc_hd__a21bo_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21bo_2

.SUBCKT sky130_fd_sc_hd__a2bb2o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a2bb2o_2

.SUBCKT sky130_fd_sc_hd__a22oi_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22oi_2

.SUBCKT sky130_fd_sc_hd__a311o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a311o_2

.SUBCKT sky130_fd_sc_hd__a21oi_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21oi_2

.SUBCKT sky130_fd_sc_hd__a21o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__a21o_2

.SUBCKT sky130_fd_sc_hd__o221a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o221a_2

.SUBCKT sky130_fd_sc_hd__conb_1 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__conb_1

.SUBCKT sky130_fd_sc_hd__einvp_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__einvp_1

.SUBCKT sky130_fd_sc_hd__o21a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21a_2

.SUBCKT sky130_fd_sc_hd__or3_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__or3_2

.SUBCKT sky130_fd_sc_hd__decap_8 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_8

.SUBCKT sky130_fd_sc_hd__or4_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__or4_2

.SUBCKT sky130_fd_sc_hd__clkbuf_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_2

.SUBCKT sky130_fd_sc_hd__nand2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nand2_2

.SUBCKT sky130_fd_sc_hd__and2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__and2_2

.SUBCKT sky130_fd_sc_hd__einvp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__einvp_2

.SUBCKT sky130_fd_sc_hd__o311a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o311a_2

.SUBCKT sky130_fd_sc_hd__and3_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__and3_2

.SUBCKT sky130_fd_sc_hd__einvn_4 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__einvn_4

.SUBCKT sky130_fd_sc_hd__einvn_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__einvn_8

.SUBCKT sky130_fd_sc_hd__o31a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o31a_2

.SUBCKT sky130_fd_sc_hd__o41a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o41a_2

.SUBCKT sky130_fd_sc_hd__decap_4 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_4

.SUBCKT sky130_fd_sc_hd__a31o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a31o_2

.SUBCKT sky130_fd_sc_hd__inv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__inv_2

.SUBCKT sky130_fd_sc_hd__mux2_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__mux2_1

.SUBCKT sky130_fd_sc_hd__o32a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__o32a_2

.SUBCKT sky130_fd_sc_hd__a32o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a32o_2

.SUBCKT sky130_fd_sc_hd__clkbuf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkbuf_1

.SUBCKT sky130_fd_sc_hd__o21ai_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__o21ai_2

.SUBCKT sky130_fd_sc_hd__tapvpwrvgnd_1 nc_1 nc_2
.ENDS sky130_fd_sc_hd__tapvpwrvgnd_1

.SUBCKT sky130_fd_sc_hd__decap_6 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_6

.SUBCKT sky130_fd_sc_hd__nor2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__nor2_2

.SUBCKT sky130_fd_sc_hd__decap_12 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_12

.SUBCKT sky130_fd_sc_hd__fill_2 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_2

.SUBCKT sky130_fd_sc_hd__diode_2 nc_1 nc_2 nc_3 nc_4 nc_5
.ENDS sky130_fd_sc_hd__diode_2

.SUBCKT sky130_fd_sc_hd__clkinv_8 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_8

.SUBCKT sky130_fd_sc_hd__clkinv_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_2

.SUBCKT sky130_fd_sc_hd__clkinv_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__clkinv_1

.SUBCKT sky130_fd_sc_hd__decap_3 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__decap_3

.SUBCKT sky130_fd_sc_hd__a221o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
+ nc_10
.ENDS sky130_fd_sc_hd__a221o_2

.SUBCKT sky130_fd_sc_hd__or2_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7
.ENDS sky130_fd_sc_hd__or2_2

.SUBCKT sky130_fd_sc_hd__fill_1 nc_1 nc_2 nc_3 nc_4
.ENDS sky130_fd_sc_hd__fill_1

.SUBCKT sky130_fd_sc_hd__a22o_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__a22o_2

.SUBCKT sky130_fd_sc_hd__o2bb2a_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8 nc_9
.ENDS sky130_fd_sc_hd__o2bb2a_2

.SUBCKT sky130_fd_sc_hd__buf_1 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6
.ENDS sky130_fd_sc_hd__buf_1

.SUBCKT sky130_fd_sc_hd__dfrtp_2 nc_1 nc_2 nc_3 nc_4 nc_5 nc_6 nc_7 nc_8
.ENDS sky130_fd_sc_hd__dfrtp_2
