*SPICE netlist created from verilog structural netlist module caravel_clocking by vlog2Spice (qflow)
*This file may contain array delimiters, not for use in simulation.

.include /home/marwan/klayout_lvs/lvs/test_cases/caravel_clocking/sky130_fd_sc_hd.spice

.subckt caravel_clocking VGND VPWR core_clk ext_clk ext_clk_sel ext_reset pll_clk
+ pll_clk90 resetb resetb_sync user_clk sel[0] sel[1] sel[2] sel2[0]
+ sel2[1] sel2[2] 

XANTENNA__283__A2 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__322__A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__323__B_N net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__347__S net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__349__B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__421__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__422__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__425__A1 net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__439__D net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__445__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__446__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__447__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__448__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__449__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__450__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__451__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__452__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__453__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__454__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__455__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__456__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__457__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__458__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__459__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__460__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__461__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__462__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__463__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__464__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__465__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__466__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__467__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__468__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__469__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__470__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__471__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__472__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__473__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__474__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__475__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__476__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__477__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__478__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__479__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__480__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__481__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__482__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__483__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__484__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__485__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__486__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__487__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__488__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__489__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__490__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__491__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__492__SET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__493__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__494__RESET_B net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_ext_clk_A ext_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_pll_clk90_A pll_clk90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_0_pll_clk_A pll_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input1_A ext_clk_sel VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input2_A ext_reset VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input3_A resetb VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input4_A sel2[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input5_A sel2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input6_A sel2[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input7_A sel[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input8_A sel[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_input9_A sel[2] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_216_ _016_ \divider2.even_0.counter[1]\ \divider2.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _121_ sky130_fd_sc_hd__mux2_1
X_217_ _121_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__clkbuf_1
X_218_ _015_ \divider2.even_0.counter[0]\ \divider2.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _122_ sky130_fd_sc_hd__mux2_1
X_219_ _122_ VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__clkbuf_1
X_220_ \divider2.even_0.N[1]\ \divider2.odd_0.old_N[1]\ VGND VGND VPWR VPWR 
+ _123_
+ sky130_fd_sc_hd__or2b_1
X_221_ \divider2.odd_0.old_N[1]\ \divider2.even_0.N[1]\ VGND VGND VPWR VPWR 
+ _124_
+ sky130_fd_sc_hd__or2b_1
X_222_ _123_ _124_ \divider2.odd_0.old_N[0]\ VGND VGND VPWR 
+ VPWR
+ _125_ sky130_fd_sc_hd__nand3_1
X_223_ \divider2.even_0.N[2]\ \divider2.odd_0.old_N[2]\ VGND VGND VPWR VPWR 
+ _126_
+ sky130_fd_sc_hd__nor2_1
X_224_ \divider2.even_0.N[2]\ \divider2.odd_0.old_N[2]\ VGND VGND VPWR VPWR 
+ _127_
+ sky130_fd_sc_hd__and2_1
X_225_ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ \divider2.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _128_ sky130_fd_sc_hd__o21a_1
X_226_ _126_ _127_ _128_ VGND VGND VPWR 
+ VPWR
+ _129_ sky130_fd_sc_hd__o21ai_1
X_227_ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ \divider2.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _130_ sky130_fd_sc_hd__o21ai_1
X_228_ \divider2.odd_0.rst_pulse\ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__clkinv_4
X_229_ _130_ _131_ VGND VGND VPWR VPWR 
+ _000_
+ sky130_fd_sc_hd__nand2_2
X_230_ _125_ _129_ _000_ VGND VGND VPWR 
+ VPWR
+ _117_ sky130_fd_sc_hd__o21a_1
X_231_ \divider2.odd_0.counter[2]\ \divider2.odd_0.counter[1]\ VGND VGND VPWR VPWR 
+ _132_
+ sky130_fd_sc_hd__nor2_1
X_232_ _132_ \divider2.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _133_
+ sky130_fd_sc_hd__nand2_1
X_233_ \divider2.odd_0.out_counter\ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__inv_2
X_234_ _133_ _134_ _128_ VGND VGND VPWR 
+ VPWR
+ _135_ sky130_fd_sc_hd__nand3b_1
X_235_ _131_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__clkbuf_2
X_236_ _130_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__clkbuf_2
X_237_ _137_ _133_ _134_ VGND VGND VPWR 
+ VPWR
+ _138_ sky130_fd_sc_hd__o21bai_1
X_238_ _135_ _136_ _138_ VGND VGND VPWR 
+ VPWR
+ _116_ sky130_fd_sc_hd__nand3_1
X_239_ _137_ _136_ \divider2.odd_0.counter[2]\ VGND VGND VPWR 
+ VPWR
+ _139_ sky130_fd_sc_hd__nand3_1
X_240_ _022_ _000_ _139_ VGND VGND VPWR 
+ VPWR
+ _115_ sky130_fd_sc_hd__a21bo_1
X_241_ _137_ _131_ \divider2.odd_0.counter[1]\ VGND VGND VPWR 
+ VPWR
+ _140_ sky130_fd_sc_hd__nand3_1
X_242_ _021_ _000_ _140_ VGND VGND VPWR 
+ VPWR
+ _114_ sky130_fd_sc_hd__a21bo_1
X_243_ _137_ _131_ \divider2.odd_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _141_ sky130_fd_sc_hd__nand3_1
X_244_ _020_ _000_ _141_ VGND VGND VPWR 
+ VPWR
+ _113_ sky130_fd_sc_hd__a21bo_1
X_245_ \divider2.odd_0.initial_begin[2]\ _025_ _002_ VGND VGND VPWR 
+ VPWR
+ _142_ sky130_fd_sc_hd__mux2_1
X_246_ _142_ VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__clkbuf_1
X_247__1 clknet_1_0_0_pll_clk90 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__inv_4
X_248_ \divider2.odd_0.initial_begin[1]\ _024_ _002_ VGND VGND VPWR 
+ VPWR
+ _143_ sky130_fd_sc_hd__mux2_1
X_249_ _143_ VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__clkbuf_1
X_250_ \divider2.odd_0.initial_begin[0]\ _023_ _002_ VGND VGND VPWR 
+ VPWR
+ _144_ sky130_fd_sc_hd__mux2_1
X_251_ _144_ VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__clkbuf_1
X_252__2 clknet_1_0_0_pll_clk90 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__inv_4
X_253_ \divider2.odd_0.initial_begin[2]\ \divider2.odd_0.initial_begin[1]\ VGND VGND VPWR VPWR 
+ _145_
+ sky130_fd_sc_hd__nor2_1
X_254_ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ \divider2.even_0.N[0]\ _145_ VGND VGND 
+ VPWR
+ VPWR _033_ sky130_fd_sc_hd__o211a_1
X_255_ \divider2.odd_0.out_counter2\ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__inv_2
X_256_ \divider2.odd_0.counter2[2]\ \divider2.odd_0.counter2[1]\ \divider2.odd_0.counter2[0]\ VGND VGND VPWR 
+ VPWR
+ _034_ sky130_fd_sc_hd__nor3b_2
X_257_ _033_ _146_ _034_ VGND VGND VPWR 
+ VPWR
+ _147_ sky130_fd_sc_hd__nand3_1
X_258_ \divider2.odd_0.counter2[2]\ \divider2.odd_0.counter2[1]\ VGND VGND VPWR VPWR 
+ _148_
+ sky130_fd_sc_hd__nor2_1
X_259_ _148_ \divider2.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _149_
+ sky130_fd_sc_hd__nand2_1
X_260_ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ \divider2.even_0.N[0]\ _145_ VGND VGND 
+ VPWR
+ VPWR _150_ sky130_fd_sc_hd__o211ai_4
X_261_ _149_ _150_ _146_ VGND VGND VPWR 
+ VPWR
+ _151_ sky130_fd_sc_hd__o21bai_1
X_262_ _147_ _151_ _136_ VGND VGND VPWR 
+ VPWR
+ _109_ sky130_fd_sc_hd__nand3_1
X_263_ _150_ _131_ VGND VGND VPWR VPWR 
+ _152_
+ sky130_fd_sc_hd__nand2_1
X_264_ _152_ _019_ VGND VGND VPWR VPWR 
+ _153_
+ sky130_fd_sc_hd__nand2_1
X_265_ _150_ _136_ \divider2.odd_0.counter2[2]\ VGND VGND VPWR 
+ VPWR
+ _154_ sky130_fd_sc_hd__nand3_1
X_266_ _153_ _154_ VGND VGND VPWR VPWR 
+ _108_
+ sky130_fd_sc_hd__nand2_1
X_267__3 clknet_1_0_0_pll_clk90 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__inv_4
X_268_ _152_ _018_ VGND VGND VPWR VPWR 
+ _155_
+ sky130_fd_sc_hd__nand2_1
X_269_ _150_ _136_ \divider2.odd_0.counter2[1]\ VGND VGND VPWR 
+ VPWR
+ _156_ sky130_fd_sc_hd__nand3_1
X_270_ _155_ _156_ VGND VGND VPWR VPWR 
+ _107_
+ sky130_fd_sc_hd__nand2_1
X_271_ \divider2.odd_0.counter2[0]\ VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__inv_2
X_272_ _152_ _017_ VGND VGND VPWR VPWR 
+ _157_
+ sky130_fd_sc_hd__nand2_1
X_273_ _065_ _152_ _157_ VGND VGND VPWR 
+ VPWR
+ _106_ sky130_fd_sc_hd__o21ai_1
X_274_ \divider2.even_0.counter[1]\ \divider2.even_0.counter[2]\ \divider2.even_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _032_ sky130_fd_sc_hd__nor3b_2
X_275_ \divider2.even_0.N[0]\ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__clkinv_4
X_276_ \divider2.even_0.out_counter\ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__clkinv_4
X_277_ _032_ _158_ _159_ VGND VGND VPWR 
+ VPWR
+ _160_ sky130_fd_sc_hd__a21o_1
X_278_ _032_ _158_ _159_ VGND VGND VPWR 
+ VPWR
+ _161_ sky130_fd_sc_hd__nand3_1
X_279_ _160_ _161_ VGND VGND VPWR VPWR 
+ _105_
+ sky130_fd_sc_hd__nand2_1
X_280_ \divider.odd_0.counter[2]\ \divider.odd_0.counter[1]\ VGND VGND VPWR VPWR 
+ _162_
+ sky130_fd_sc_hd__nor2_1
X_281_ _162_ \divider.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _163_
+ sky130_fd_sc_hd__nand2_1
X_282_ \divider.odd_0.out_counter\ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__inv_2
X_283_ net30 net26 \divider.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _165_ sky130_fd_sc_hd__o21a_1
X_284_ _163_ _164_ _165_ VGND VGND VPWR 
+ VPWR
+ _166_ sky130_fd_sc_hd__nand3b_1
X_285_ \divider.odd_0.rst_pulse\ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__clkinv_4
X_286_ _167_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__clkbuf_2
X_287_ \divider.even_0.N[2]\ \divider.even_0.N[1]\ \divider.even_0.N[0]\ VGND VGND VPWR 
+ VPWR
+ _169_ sky130_fd_sc_hd__o21ai_1
X_288_ _169_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__clkbuf_2
X_289_ _170_ _163_ _164_ VGND VGND VPWR 
+ VPWR
+ _171_ sky130_fd_sc_hd__o21bai_1
X_290_ _166_ _168_ _171_ VGND VGND VPWR 
+ VPWR
+ _104_ sky130_fd_sc_hd__nand3_1
X_291_ _169_ _167_ VGND VGND VPWR VPWR 
+ _001_
+ sky130_fd_sc_hd__nand2_2
X_292_ _170_ \divider.odd_0.counter[2]\ _168_ VGND VGND VPWR 
+ VPWR
+ _172_ sky130_fd_sc_hd__nand3_1
X_293_ _011_ _001_ _172_ VGND VGND VPWR 
+ VPWR
+ _103_ sky130_fd_sc_hd__a21bo_1
X_294_ _170_ \divider.odd_0.counter[1]\ _167_ VGND VGND VPWR 
+ VPWR
+ _173_ sky130_fd_sc_hd__nand3_1
X_295_ _010_ _001_ _173_ VGND VGND VPWR 
+ VPWR
+ _102_ sky130_fd_sc_hd__a21bo_1
X_296_ _170_ \divider.odd_0.counter[0]\ _167_ VGND VGND VPWR 
+ VPWR
+ _174_ sky130_fd_sc_hd__nand3_1
X_297_ _009_ _001_ _174_ VGND VGND VPWR 
+ VPWR
+ _101_ sky130_fd_sc_hd__a21bo_1
X_298_ \divider.odd_0.initial_begin[2]\ _014_ _003_ VGND VGND VPWR 
+ VPWR
+ _175_ sky130_fd_sc_hd__mux2_1
X_299_ _175_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__clkbuf_1
X_300__4 clknet_1_0_0_pll_clk VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__inv_4
X_301_ \divider.odd_0.initial_begin[1]\ _013_ _003_ VGND VGND VPWR 
+ VPWR
+ _176_ sky130_fd_sc_hd__mux2_1
X_302_ _176_ VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__clkbuf_1
X_303_ \divider.odd_0.initial_begin[0]\ _012_ _003_ VGND VGND VPWR 
+ VPWR
+ _177_ sky130_fd_sc_hd__mux2_1
X_304_ _177_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__clkbuf_1
X_305__5 clknet_1_1_0_pll_clk VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__inv_4
X_306_ \divider.odd_0.initial_begin[2]\ \divider.odd_0.initial_begin[1]\ VGND VGND VPWR VPWR 
+ _178_
+ sky130_fd_sc_hd__nor2_1
X_307_ \divider.even_0.N[2]\ \divider.even_0.N[1]\ \divider.even_0.N[0]\ _178_ VGND VGND 
+ VPWR
+ VPWR _029_ sky130_fd_sc_hd__o211a_1
X_308_ \divider.odd_0.out_counter2\ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__inv_2
X_309_ \divider.odd_0.counter2[2]\ \divider.odd_0.counter2[1]\ \divider.odd_0.counter2[0]\ VGND VGND VPWR 
+ VPWR
+ _030_ sky130_fd_sc_hd__nor3b_2
X_310_ net38 _179_ _030_ VGND VGND VPWR 
+ VPWR
+ _180_ sky130_fd_sc_hd__nand3_1
X_311_ \divider.odd_0.counter2[2]\ \divider.odd_0.counter2[1]\ VGND VGND VPWR VPWR 
+ _181_
+ sky130_fd_sc_hd__nor2_1
X_312_ _181_ \divider.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _182_
+ sky130_fd_sc_hd__nand2_1
X_313_ net27 net28 net32 _178_ VGND VGND 
+ VPWR
+ VPWR _183_ sky130_fd_sc_hd__o211ai_4
X_314_ _182_ _183_ _179_ VGND VGND VPWR 
+ VPWR
+ _184_ sky130_fd_sc_hd__o21bai_1
X_315_ _180_ _184_ _168_ VGND VGND VPWR 
+ VPWR
+ _097_ sky130_fd_sc_hd__nand3_1
X_316_ \divider.even_0.N[0]\ \divider.even_0.counter[1]\ \divider.even_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _185_ sky130_fd_sc_hd__nor3_1
X_317_ \divider.even_0.counter[2]\ _185_ VGND VGND VPWR VPWR 
+ _096_
+ sky130_fd_sc_hd__xor2_1
X_318_ _005_ \divider.even_0.counter[1]\ net34 VGND VGND VPWR 
+ VPWR
+ _186_ sky130_fd_sc_hd__mux2_1
X_319_ _186_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__clkbuf_1
X_320_ _004_ \divider.even_0.counter[0]\ net34 VGND VGND VPWR 
+ VPWR
+ _187_ sky130_fd_sc_hd__mux2_1
X_321_ _187_ VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__clkbuf_1
X_322_ net26 \divider.odd_0.old_N[1]\ VGND VGND VPWR VPWR 
+ _188_
+ sky130_fd_sc_hd__or2b_1
X_323_ \divider.odd_0.old_N[1]\ net26 VGND VGND VPWR VPWR 
+ _189_
+ sky130_fd_sc_hd__or2b_1
X_324_ _188_ _189_ \divider.odd_0.old_N[0]\ VGND VGND VPWR 
+ VPWR
+ _190_ sky130_fd_sc_hd__nand3_1
X_325_ net30 \divider.odd_0.old_N[2]\ VGND VGND VPWR VPWR 
+ _191_
+ sky130_fd_sc_hd__nor2_1
X_326_ net30 \divider.odd_0.old_N[2]\ VGND VGND VPWR VPWR 
+ _192_
+ sky130_fd_sc_hd__and2_1
X_327_ _191_ _192_ _165_ VGND VGND VPWR 
+ VPWR
+ _193_ sky130_fd_sc_hd__o21ai_1
X_328_ _190_ _193_ _001_ VGND VGND VPWR 
+ VPWR
+ _093_ sky130_fd_sc_hd__o21a_1
X_329_ _183_ _167_ VGND VGND VPWR VPWR 
+ _194_
+ sky130_fd_sc_hd__nand2_1
X_330_ _194_ _008_ VGND VGND VPWR VPWR 
+ _195_
+ sky130_fd_sc_hd__nand2_1
X_331_ _183_ _168_ \divider.odd_0.counter2[2]\ VGND VGND VPWR 
+ VPWR
+ _196_ sky130_fd_sc_hd__nand3_1
X_332_ _195_ _196_ VGND VGND VPWR VPWR 
+ _092_
+ sky130_fd_sc_hd__nand2_1
X_333__6 clknet_1_1_0_pll_clk VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__inv_4
X_334_ _194_ _007_ VGND VGND VPWR VPWR 
+ _197_
+ sky130_fd_sc_hd__nand2_1
X_335_ _183_ _168_ \divider.odd_0.counter2[1]\ VGND VGND VPWR 
+ VPWR
+ _198_ sky130_fd_sc_hd__nand3_1
X_336_ _197_ _198_ VGND VGND VPWR VPWR 
+ _091_
+ sky130_fd_sc_hd__nand2_1
X_337_ \divider.odd_0.counter2[0]\ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__inv_2
X_338_ _194_ _006_ VGND VGND VPWR VPWR 
+ _199_
+ sky130_fd_sc_hd__nand2_1
X_339_ _045_ _194_ _199_ VGND VGND VPWR 
+ VPWR
+ _090_ sky130_fd_sc_hd__o21ai_1
X_340_ \divider.even_0.counter[2]\ \divider.even_0.counter[1]\ VGND VGND VPWR VPWR 
+ _200_
+ sky130_fd_sc_hd__nor2_1
X_341_ net31 VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__clkinv_4
X_342_ _200_ _201_ \divider.even_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _202_ sky130_fd_sc_hd__nand3_1
X_343_ \divider.even_0.out_counter\ _202_ VGND VGND VPWR VPWR 
+ _089_
+ sky130_fd_sc_hd__xnor2_1
X_344__9 net10 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__inv_4
X_345__8 net10 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__inv_4
X_346__7 net10 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__inv_4
X_347_ ext_clk_syncd_pre clknet_1_0_0_ext_clk net3 VGND VGND VPWR 
+ VPWR
+ _203_ sky130_fd_sc_hd__mux2_2
X_348_ _203_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__buf_1
X_349_ net30 net26 VGND VGND VPWR VPWR 
+ _026_
+ sky130_fd_sc_hd__nor2_1
X_350_ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ VGND VGND VPWR VPWR 
+ _027_
+ sky130_fd_sc_hd__nor2_1
X_351_ \divider.even_0.counter[2]\ \divider.even_0.counter[1]\ \divider.even_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _028_ sky130_fd_sc_hd__nor3b_1
X_352_ _163_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkinv_4
X_353_ _133_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkinv_4
X_354_ \divider.odd_0.out_counter\ \divider.odd_0.out_counter2\ VGND VGND VPWR VPWR 
+ _204_
+ sky130_fd_sc_hd__xnor2_1
X_355_ _201_ _036_ _170_ _204_ VGND VGND 
+ VPWR
+ VPWR \divider.out\ sky130_fd_sc_hd__o2bb2ai_2
X_356_ \divider2.odd_0.out_counter\ \divider2.odd_0.out_counter2\ VGND VGND VPWR VPWR 
+ _205_
+ sky130_fd_sc_hd__xnor2_1
X_357_ _158_ _038_ _137_ _205_ VGND VGND 
+ VPWR
+ VPWR \divider2.out\ sky130_fd_sc_hd__o2bb2ai_2
X_358_ \divider.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__clkinv_2
X_359_ net33 net29 VGND VGND VPWR VPWR 
+ _040_
+ sky130_fd_sc_hd__xnor2_1
X_360_ \divider.odd_0.initial_begin[1]\ \divider.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR 
+ _041_
+ sky130_fd_sc_hd__xnor2_1
X_361_ net33 \divider.even_0.N[2]\ net29 VGND VGND VPWR 
+ VPWR
+ _206_ sky130_fd_sc_hd__nor3_1
X_362_ net33 net29 \divider.even_0.N[2]\ VGND VGND VPWR 
+ VPWR
+ _044_ sky130_fd_sc_hd__o21a_1
X_363_ _206_ _044_ VGND VGND VPWR VPWR 
+ _042_
+ sky130_fd_sc_hd__nor2_1
X_364_ \divider.odd_0.initial_begin[1]\ \divider.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR 
+ _207_
+ sky130_fd_sc_hd__nor2_1
X_365_ \divider.odd_0.initial_begin[2]\ _207_ VGND VGND VPWR VPWR 
+ _043_
+ sky130_fd_sc_hd__xor2_1
X_366_ \divider.odd_0.counter2[1]\ \divider.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _047_
+ sky130_fd_sc_hd__xnor2_1
X_367_ \divider.odd_0.counter2[1]\ \divider.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _208_
+ sky130_fd_sc_hd__nor2_1
X_368_ \divider.odd_0.counter2[2]\ _208_ VGND VGND VPWR VPWR 
+ _049_
+ sky130_fd_sc_hd__xor2_1
X_369_ \divider.odd_0.counter[0]\ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkinv_2
X_370_ \divider.odd_0.counter[1]\ \divider.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _053_
+ sky130_fd_sc_hd__xnor2_1
X_371_ \divider.odd_0.counter[1]\ \divider.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _209_
+ sky130_fd_sc_hd__nor2_1
X_372_ \divider.odd_0.counter[2]\ _209_ VGND VGND VPWR VPWR 
+ _055_
+ sky130_fd_sc_hd__xor2_1
X_373_ \divider.even_0.counter[0]\ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__clkinv_2
X_374_ \divider.even_0.counter[1]\ \divider.even_0.counter[0]\ VGND VGND VPWR VPWR 
+ _058_
+ sky130_fd_sc_hd__xnor2_1
X_375_ \divider2.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__clkinv_2
X_376_ \divider2.even_0.N[0]\ \divider2.even_0.N[1]\ VGND VGND VPWR VPWR 
+ _060_
+ sky130_fd_sc_hd__xnor2_1
X_377_ \divider2.odd_0.initial_begin[1]\ \divider2.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR 
+ _061_
+ sky130_fd_sc_hd__xnor2_1
X_378_ \divider2.even_0.N[0]\ \divider2.even_0.N[2]\ \divider2.even_0.N[1]\ VGND VGND VPWR 
+ VPWR
+ _210_ sky130_fd_sc_hd__nor3_1
X_379_ \divider2.even_0.N[0]\ \divider2.even_0.N[1]\ \divider2.even_0.N[2]\ VGND VGND VPWR 
+ VPWR
+ _064_ sky130_fd_sc_hd__o21a_1
X_380_ _210_ _064_ VGND VGND VPWR VPWR 
+ _062_
+ sky130_fd_sc_hd__nor2_1
X_381_ \divider2.odd_0.initial_begin[1]\ \divider2.odd_0.initial_begin[0]\ VGND VGND VPWR VPWR 
+ _211_
+ sky130_fd_sc_hd__nor2_1
X_382_ \divider2.odd_0.initial_begin[2]\ _211_ VGND VGND VPWR VPWR 
+ _063_
+ sky130_fd_sc_hd__xor2_1
X_383_ \divider2.odd_0.counter2[1]\ \divider2.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _067_
+ sky130_fd_sc_hd__xnor2_1
X_384_ \divider2.odd_0.counter2[1]\ \divider2.odd_0.counter2[0]\ VGND VGND VPWR VPWR 
+ _212_
+ sky130_fd_sc_hd__nor2_1
X_385_ \divider2.odd_0.counter2[2]\ _212_ VGND VGND VPWR VPWR 
+ _069_
+ sky130_fd_sc_hd__xor2_1
X_386_ \divider2.odd_0.counter[0]\ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__clkinv_2
X_387_ \divider2.odd_0.counter[1]\ \divider2.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _073_
+ sky130_fd_sc_hd__xnor2_1
X_388_ \divider2.odd_0.counter[1]\ \divider2.odd_0.counter[0]\ VGND VGND VPWR VPWR 
+ _213_
+ sky130_fd_sc_hd__nor2_1
X_389_ \divider2.odd_0.counter[2]\ _213_ VGND VGND VPWR VPWR 
+ _075_
+ sky130_fd_sc_hd__xor2_1
X_390_ \divider2.even_0.counter[0]\ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__clkinv_2
X_391_ \divider2.even_0.counter[1]\ \divider2.even_0.counter[0]\ VGND VGND VPWR VPWR 
+ _078_
+ sky130_fd_sc_hd__xnor2_1
X_392_ net1 VGND VGND VPWR VPWR pll_clk_sel sky130_fd_sc_hd__clkinv_4
X_393_ net2 \reset_delay[0]\ VGND VGND VPWR VPWR 
+ net11
+ sky130_fd_sc_hd__nor2_1
X_394_ \divider2.even_0.counter[1]\ \divider2.even_0.N[0]\ \divider2.even_0.counter[0]\ VGND VGND VPWR 
+ VPWR
+ _214_ sky130_fd_sc_hd__nor3_1
X_395_ \divider2.even_0.counter[2]\ _214_ VGND VGND VPWR VPWR 
+ _120_
+ sky130_fd_sc_hd__xor2_1
X_396__13 VGND VGND VPWR VPWR NC net13 sky130_fd_sc_hd__conb_1
X_397_ _000_ \divider2.odd_0.rst_pulse\ _033_ VGND VGND VPWR 
+ VPWR
+ _002_ sky130_fd_sc_hd__mux2_1
X_398_ _001_ \divider.odd_0.rst_pulse\ _029_ VGND VGND VPWR 
+ VPWR
+ _003_ sky130_fd_sc_hd__mux2_2
X_399_ _037_ \divider.out\ use_pll_second VGND VGND VPWR 
+ VPWR
+ net10 sky130_fd_sc_hd__mux2_1
X_400_ _037_ \divider2.out\ use_pll_second VGND VGND VPWR 
+ VPWR
+ net12 sky130_fd_sc_hd__mux2_1
X_401_ _065_ \divider2.even_0.N[0]\ _034_ VGND VGND VPWR 
+ VPWR
+ _066_ sky130_fd_sc_hd__mux2_1
X_402_ _066_ \divider2.even_0.N[0]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _017_ sky130_fd_sc_hd__mux2_1
X_403_ _067_ \divider2.even_0.N[1]\ _034_ VGND VGND VPWR 
+ VPWR
+ _068_ sky130_fd_sc_hd__mux2_1
X_404_ _068_ \divider2.even_0.N[1]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _018_ sky130_fd_sc_hd__mux2_1
X_405_ _073_ \divider2.even_0.N[1]\ _035_ VGND VGND VPWR 
+ VPWR
+ _074_ sky130_fd_sc_hd__mux2_1
X_406_ _074_ \divider2.even_0.N[1]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _021_ sky130_fd_sc_hd__mux2_1
X_407_ _075_ \divider2.even_0.N[2]\ _035_ VGND VGND VPWR 
+ VPWR
+ _076_ sky130_fd_sc_hd__mux2_1
X_408_ _076_ \divider2.even_0.N[2]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _022_ sky130_fd_sc_hd__mux2_1
X_409_ _077_ \divider2.even_0.N[1]\ _032_ VGND VGND VPWR 
+ VPWR
+ _015_ sky130_fd_sc_hd__mux2_1
X_410_ _039_ _040_ \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _012_ sky130_fd_sc_hd__mux2_1
X_411_ _041_ _042_ \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _013_ sky130_fd_sc_hd__mux2_1
X_412_ _043_ _044_ \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _014_ sky130_fd_sc_hd__mux2_1
X_413_ _045_ \divider.even_0.N[0]\ _030_ VGND VGND VPWR 
+ VPWR
+ _046_ sky130_fd_sc_hd__mux2_1
X_414_ _046_ \divider.even_0.N[0]\ \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _006_ sky130_fd_sc_hd__mux2_1
X_415_ _047_ \divider.even_0.N[1]\ _030_ VGND VGND VPWR 
+ VPWR
+ _048_ sky130_fd_sc_hd__mux2_1
X_416_ _048_ \divider.even_0.N[1]\ \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _007_ sky130_fd_sc_hd__mux2_1
X_417_ _049_ \divider.even_0.N[2]\ _030_ VGND VGND VPWR 
+ VPWR
+ _050_ sky130_fd_sc_hd__mux2_1
X_418_ _050_ net37 \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _008_ sky130_fd_sc_hd__mux2_1
X_419_ _051_ net35 _031_ VGND VGND VPWR 
+ VPWR
+ _052_ sky130_fd_sc_hd__mux2_1
X_420_ _052_ net36 \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _009_ sky130_fd_sc_hd__mux2_1
X_421_ _053_ net26 _031_ VGND VGND VPWR 
+ VPWR
+ _054_ sky130_fd_sc_hd__mux2_1
X_422_ _054_ net26 \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _010_ sky130_fd_sc_hd__mux2_1
X_423_ _055_ net37 _031_ VGND VGND VPWR 
+ VPWR
+ _056_ sky130_fd_sc_hd__mux2_1
X_424_ _056_ net30 \divider.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _011_ sky130_fd_sc_hd__mux2_1
X_425_ _057_ net26 _028_ VGND VGND VPWR 
+ VPWR
+ _004_ sky130_fd_sc_hd__mux2_1
X_426_ _058_ net30 _028_ VGND VGND VPWR 
+ VPWR
+ _005_ sky130_fd_sc_hd__mux2_1
X_427_ _059_ _060_ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _023_ sky130_fd_sc_hd__mux2_1
X_428_ _061_ _062_ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _024_ sky130_fd_sc_hd__mux2_1
X_429_ _063_ _064_ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _025_ sky130_fd_sc_hd__mux2_1
X_430_ _069_ \divider2.even_0.N[2]\ _034_ VGND VGND VPWR 
+ VPWR
+ _070_ sky130_fd_sc_hd__mux2_1
X_431_ _070_ \divider2.even_0.N[2]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _019_ sky130_fd_sc_hd__mux2_1
X_432_ _071_ \divider2.even_0.N[0]\ _035_ VGND VGND VPWR 
+ VPWR
+ _072_ sky130_fd_sc_hd__mux2_1
X_433_ _072_ \divider2.even_0.N[0]\ \divider2.odd_0.rst_pulse\ VGND VGND VPWR 
+ VPWR
+ _020_ sky130_fd_sc_hd__mux2_1
X_434_ _078_ \divider2.even_0.N[2]\ _032_ VGND VGND VPWR 
+ VPWR
+ _016_ sky130_fd_sc_hd__mux2_1
X_435_ \divider.even_0.out_counter\ clknet_1_1_0_pll_clk _026_ VGND VGND VPWR 
+ VPWR
+ _036_ sky130_fd_sc_hd__mux2_1
X_436_ clknet_1_1_0_ext_clk ext_clk_syncd use_pll_first VGND VGND VPWR 
+ VPWR
+ _037_ sky130_fd_sc_hd__mux2_1
X_437_ \divider2.even_0.out_counter\ clknet_1_1_0_pll_clk90 _027_ VGND VGND VPWR 
+ VPWR
+ _038_ sky130_fd_sc_hd__mux2_1
X_438_ clknet_1_1_0_pll_clk \divider.even_0.N[0]\ VGND VGND VPWR VPWR 
+ \divider.odd_0.old_N[0]\
+ sky130_fd_sc_hd__dfxtp_1
X_439_ clknet_1_1_0_pll_clk net26 VGND VGND VPWR VPWR 
+ \divider.odd_0.old_N[1]\
+ sky130_fd_sc_hd__dfxtp_1
X_440_ clknet_1_1_0_pll_clk net30 VGND VGND VPWR VPWR 
+ \divider.odd_0.old_N[2]\
+ sky130_fd_sc_hd__dfxtp_1
X_441_ clknet_1_1_0_pll_clk90 \divider2.even_0.N[0]\ VGND VGND VPWR VPWR 
+ \divider2.odd_0.old_N[0]\
+ sky130_fd_sc_hd__dfxtp_1
X_442_ clknet_1_0_0_pll_clk90 \divider2.even_0.N[1]\ VGND VGND VPWR VPWR 
+ \divider2.odd_0.old_N[1]\
+ sky130_fd_sc_hd__dfxtp_1
X_443_ clknet_1_1_0_pll_clk90 \divider2.even_0.N[2]\ VGND VGND VPWR VPWR 
+ \divider2.odd_0.old_N[2]\
+ sky130_fd_sc_hd__dfxtp_1
X_444_ clknet_1_0_0_pll_clk _088_ VGND VGND VPWR VPWR 
+ ext_clk_syncd_pre
+ sky130_fd_sc_hd__dfxtp_1
X_445_ net20 net25 net3 VGND VGND VPWR 
+ VPWR
+ \reset_delay[0]\ sky130_fd_sc_hd__dfstp_1
X_446_ net21 net24 net3 VGND VGND VPWR 
+ VPWR
+ \reset_delay[1]\ sky130_fd_sc_hd__dfstp_1
X_447_ net22 net13 net3 VGND VGND VPWR 
+ VPWR
+ \reset_delay[2]\ sky130_fd_sc_hd__dfstp_1
X_448_ clknet_1_1_0_pll_clk pll_clk_sel net3 VGND VGND VPWR 
+ VPWR
+ use_pll_first sky130_fd_sc_hd__dfrtp_1
X_449_ clknet_1_1_0_pll_clk use_pll_first net3 VGND VGND VPWR 
+ VPWR
+ use_pll_second sky130_fd_sc_hd__dfrtp_1
X_450_ clknet_1_1_0_pll_clk net23 net3 VGND VGND VPWR 
+ VPWR
+ ext_clk_syncd sky130_fd_sc_hd__dfrtp_1
X_451_ \divider.out\ net7 net3 VGND VGND VPWR 
+ VPWR
+ \divider.syncNp[0]\ sky130_fd_sc_hd__dfrtp_1
X_452_ \divider.out\ net8 net3 VGND VGND VPWR 
+ VPWR
+ \divider.syncNp[1]\ sky130_fd_sc_hd__dfstp_1
X_453_ \divider.out\ net9 net3 VGND VGND VPWR 
+ VPWR
+ \divider.syncNp[2]\ sky130_fd_sc_hd__dfrtp_1
X_454_ \divider.out\ \divider.syncNp[0]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.N[0]\ sky130_fd_sc_hd__dfrtp_4
X_455_ \divider.out\ \divider.syncNp[1]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.N[1]\ sky130_fd_sc_hd__dfstp_4
X_456_ \divider.out\ \divider.syncNp[2]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.N[2]\ sky130_fd_sc_hd__dfrtp_4
X_457_ \divider2.out\ net4 net3 VGND VGND VPWR 
+ VPWR
+ \divider2.syncNp[0]\ sky130_fd_sc_hd__dfrtp_1
X_458_ \divider2.out\ net5 net3 VGND VGND VPWR 
+ VPWR
+ \divider2.syncNp[1]\ sky130_fd_sc_hd__dfstp_1
X_459_ \divider2.out\ net6 net3 VGND VGND VPWR 
+ VPWR
+ \divider2.syncNp[2]\ sky130_fd_sc_hd__dfrtp_1
X_460_ \divider2.out\ \divider2.syncNp[0]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.N[0]\ sky130_fd_sc_hd__dfrtp_4
X_461_ \divider2.out\ \divider2.syncNp[1]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.N[1]\ sky130_fd_sc_hd__dfstp_4
X_462_ \divider2.out\ \divider2.syncNp[2]\ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.N[2]\ sky130_fd_sc_hd__dfrtp_4
X_463_ clknet_1_1_0_pll_clk _089_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.out_counter\ sky130_fd_sc_hd__dfstp_1
X_464_ clknet_1_1_0_pll_clk _090_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter2[0]\ sky130_fd_sc_hd__dfrtn_1
X_465_ net19 _091_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter2[1]\ sky130_fd_sc_hd__dfstp_1
X_466_ clknet_1_1_0_pll_clk _092_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter2[2]\ sky130_fd_sc_hd__dfrtn_1
X_467_ clknet_1_1_0_pll_clk _093_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.rst_pulse\ sky130_fd_sc_hd__dfrtp_4
X_468_ clknet_1_0_0_pll_clk _094_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.counter[0]\ sky130_fd_sc_hd__dfstp_2
X_469_ clknet_1_0_0_pll_clk _095_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.counter[1]\ sky130_fd_sc_hd__dfrtp_2
X_470_ clknet_1_0_0_pll_clk _096_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.even_0.counter[2]\ sky130_fd_sc_hd__dfrtp_1
X_471_ net18 _097_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.out_counter2\ sky130_fd_sc_hd__dfstp_1
X_472_ clknet_1_0_0_pll_clk _098_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.initial_begin[0]\ sky130_fd_sc_hd__dfrtn_1
X_473_ net17 _099_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.initial_begin[1]\ sky130_fd_sc_hd__dfstp_1
X_474_ clknet_1_0_0_pll_clk _100_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.initial_begin[2]\ sky130_fd_sc_hd__dfrtn_1
X_475_ clknet_1_1_0_pll_clk _101_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter[0]\ sky130_fd_sc_hd__dfrtp_2
X_476_ clknet_1_0_0_pll_clk _102_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter[1]\ sky130_fd_sc_hd__dfstp_1
X_477_ clknet_1_0_0_pll_clk _103_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.counter[2]\ sky130_fd_sc_hd__dfrtp_1
X_478_ clknet_1_0_0_pll_clk _104_ net3 VGND VGND VPWR 
+ VPWR
+ \divider.odd_0.out_counter\ sky130_fd_sc_hd__dfstp_1
X_479_ clknet_1_1_0_pll_clk90 _105_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.out_counter\ sky130_fd_sc_hd__dfstp_1
X_480_ clknet_1_0_0_pll_clk90 _106_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter2[0]\ sky130_fd_sc_hd__dfrtn_1
X_481_ net16 _107_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter2[1]\ sky130_fd_sc_hd__dfstp_1
X_482_ clknet_1_0_0_pll_clk90 _108_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter2[2]\ sky130_fd_sc_hd__dfrtn_1
X_483_ net15 _109_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.out_counter2\ sky130_fd_sc_hd__dfstp_1
X_484_ clknet_1_0_0_pll_clk90 _110_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.initial_begin[0]\ sky130_fd_sc_hd__dfrtn_1
X_485_ net14 _111_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.initial_begin[1]\ sky130_fd_sc_hd__dfstp_1
X_486_ clknet_1_0_0_pll_clk90 _112_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.initial_begin[2]\ sky130_fd_sc_hd__dfrtn_1
X_487_ clknet_1_1_0_pll_clk90 _113_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter[0]\ sky130_fd_sc_hd__dfrtp_2
X_488_ clknet_1_0_0_pll_clk90 _114_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter[1]\ sky130_fd_sc_hd__dfstp_1
X_489_ clknet_1_0_0_pll_clk90 _115_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.counter[2]\ sky130_fd_sc_hd__dfrtp_1
X_490_ clknet_1_1_0_pll_clk90 _116_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.out_counter\ sky130_fd_sc_hd__dfstp_1
X_491_ clknet_1_1_0_pll_clk90 _117_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.odd_0.rst_pulse\ sky130_fd_sc_hd__dfrtp_4
X_492_ clknet_1_1_0_pll_clk90 _118_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.counter[0]\ sky130_fd_sc_hd__dfstp_1
X_493_ clknet_1_1_0_pll_clk90 _119_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.counter[1]\ sky130_fd_sc_hd__dfrtp_1
X_494_ clknet_1_1_0_pll_clk90 _120_ net3 VGND VGND VPWR 
+ VPWR
+ \divider2.even_0.counter[2]\ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_0_ext_clk ext_clk VGND VGND VPWR VPWR clknet_0_ext_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0_pll_clk pll_clk VGND VGND VPWR VPWR clknet_0_pll_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_0_pll_clk90 pll_clk90 VGND VGND VPWR VPWR clknet_0_pll_clk90 sky130_fd_sc_hd__clkbuf_16
Xclkbuf_1_0_0_ext_clk clknet_0_ext_clk VGND VGND VPWR VPWR clknet_1_0_0_ext_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0_pll_clk clknet_0_pll_clk VGND VGND VPWR VPWR clknet_1_0_0_pll_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_0_0_pll_clk90 clknet_0_pll_clk90 VGND VGND VPWR VPWR clknet_1_0_0_pll_clk90 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_ext_clk clknet_0_ext_clk VGND VGND VPWR VPWR clknet_1_1_0_ext_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_pll_clk clknet_0_pll_clk VGND VGND VPWR VPWR clknet_1_1_0_pll_clk sky130_fd_sc_hd__clkbuf_2
Xclkbuf_1_1_0_pll_clk90 clknet_0_pll_clk90 VGND VGND VPWR VPWR clknet_1_1_0_pll_clk90 sky130_fd_sc_hd__clkbuf_2
Xhold1 ext_clk_syncd_pre VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold2 \reset_delay[2]\ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold3 \reset_delay[1]\ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkdlybuf4s25_1
Xinput1 ext_clk_sel VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
Xinput2 ext_reset VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
Xinput3 resetb VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_12
Xinput4 sel2[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
Xinput5 sel2[1] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
Xinput6 sel2[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
Xinput7 sel[0] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
Xinput8 sel[1] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
Xinput9 sel[2] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
Xoutput10 net10 VGND VGND VPWR VPWR core_clk sky130_fd_sc_hd__clkbuf_1
Xoutput11 net11 VGND VGND VPWR VPWR resetb_sync sky130_fd_sc_hd__buf_2
Xoutput12 net12 VGND VGND VPWR VPWR user_clk sky130_fd_sc_hd__clkbuf_1
Xrebuffer10 \divider.even_0.N[0]\ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xrebuffer11 \divider.even_0.N[0]\ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xrebuffer12 net33 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer13 \divider.even_0.N[0]\ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer14 net35 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer16 _029_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer5 net37 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xrebuffer6 \divider.even_0.N[1]\ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dlygate4sd1_1
Xrebuffer7 \divider.even_0.N[1]\ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
Xrebuffer9 \divider.even_0.N[0]\ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xsplit15 \divider.even_0.N[2]\ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_2
Xsplit4 \divider.even_0.N[1]\ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_4
Xsplit8 net37 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_2

.ends
.end
